module mario_top
( 
	input [0:0]CLOCK_50,
	
	input [1:0]SW,
	input PS2_CLK,
	input PS2_DAT,

	output wire VGA_HS , VGA_VS ,
	output wire [3:0]VGA_R,VGA_G,VGA_B,
	output wire [9:0] mario_x_reg
); 

	wire [8:0] rgb_next; 
	reg  [8:0]rgb_reg; 
	wire [8:0]rgb;

	wire [9:0] pixel_x , pixel_y; 
	wire video_on , pixel_tick; 
	wire up,left,down,right,fast,jump;
	
	assign VGA_R = {rgb[8:6],1'b0};
	assign VGA_G = {rgb[5:3],1'b0};
	assign VGA_B = {rgb[2:0],1'b0};
	
	keyboard keyboard1(SW[1],PS2_CLK, PS2_DAT, up, down, left, right, fast, jump); //Keyboard driver
	
	vga_sync  vsync_unit (.clk(CLOCK_50[0]),  .reset (SW[1]), .hsync(VGA_HS),  .vsync(VGA_VS), .video_on(video_on),  .p_tick(pixel_tick), .pixel_x(pixel_x),  .pixel_y(pixel_y)); //VGA driver
	mario  mario1 (.CLOCK_50(CLOCK_50[0]), .reset(SW[1]), .pix_x(pixel_x),  .pix_y(pixel_y), 
				  .video_on(video_on), .KEY({up,down,fast,jump,left,right}), .graph_rgb(rgb_next)) ; // pixel color generation
	always @(posedge CLOCK_50) 
		if  (pixel_tick) rgb_reg <=  rgb_next ; 
	assign rgb = rgb_reg; 	
	
endmodule




module mario 
(	
	input wire [0:0]CLOCK_50,
	input wire reset,
	input wire [9:0]pix_x,pix_y,
	input wire video_on,
	input wire [5:0]KEY,

	output reg [8:0]graph_rgb

);
	localparam MAX_X = 640;
	localparam MAX_Y = 480;
        
    localparam BASE = MAX_Y - 1 - 50; //Base that mario stand on
	wire refr_tick;
	wire at_mid_next;
	reg  at_mid_reg;
	
	//Built Counter which used to generate scene for game
	reg [30:0] built_reg;
	wire [30:0] built_next;
	
//	--------------------------MARIO--------------------------------
	reg[9:0] mario_lo_size,mario_hi_size; //mario long size and mario high size
	reg shift;
	reg big;
	reg big_next;
	reg [9:0]vr; //run velocity
	reg [9:0] vr_next;
	reg [9:0]max_jump ; //high maximum that mario can jump
	reg [9:0]max_jump_next;
	reg [8:0]backgroud_rgb = 9'b000100111; //Blue color
	
	
	wire [9:0]mario_x_next,mario_y_next;
	reg [9:0]mario_x_reg,mario_y_reg;	
	wire [9:0] mario_x_l,mario_x_r,mario_y_t,mario_y_b;	
	reg [9:0]mario_del_run_next,mario_del_jump_next;
	reg [9:0]mario_del_jump_reg;
	reg [9:0]mario_del_run_reg;	

	reg Drop_next; //that cotrol the state drop of mario
	reg Drop_reg;
	reg [1:0] state_next;
	reg [1:0] state_reg;

	wire [9:0]mario_highest_next; //update the highest level mario can jump
	reg  [9:0]mario_highest_reg;
	reg [9:0] mario_base_reg;// update the base that mario can stand on
    wire [9:0]mario_base_next;
	

	
	//--------------------------GROUND--------------------------------
	localparam GROUND_Y_T = 430;
	localparam GROUND_Y_B = 480;
	wire ground_on;
	reg [8:0]ground_rgb = 9'b101001000; //Orange color
	
	//--------------------------PRINCESS---------1-----------------------------------
	localparam PRI_LO_SIZE = 148;
	localparam PRI_HI_SIZE = 190;
	reg [9:0] pri_x_reg;
	reg [9:0] pri_x_next;
	wire [9:0] pri_x_l, pri_x_r;
	wire [9:0] pri_y_t, pri_y_b; 
	wire [7:0] rom_addr_pri;
	wire [7:0] rom_col_pri;
	reg [150:0] rom_data_pri;
	wire rom_bit_pri;
	wire sq_pri_on, rd_pri_on;
	reg [8:0] pri_rgb = 9'b011000011; //Violet color
	
	always @*
	case(rom_addr_pri)
	
		8'd0 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'd1 : rom_data_pri  = 150'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'd2 : rom_data_pri  = 150'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		8'd3 : rom_data_pri =  150'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		8'd4 : rom_data_pri =   150'b010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
		8'd5 : rom_data_pri =  150'b001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
		8'd6 : rom_data_pri =  150'b001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
		8'd7 : rom_data_pri = 150'b000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
		8'd8 : rom_data_pri =  150'b000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000;
		8'd9 : rom_data_pri = 150'b000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
		8'd10 : rom_data_pri =   150'b000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000;
		8'd11 : rom_data_pri =   150'b000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000;
		8'd12 : rom_data_pri =  150'b000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
		8'd13 : rom_data_pri =  150'b000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000;
		8'd14 : rom_data_pri =  150'b000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000;
		8'd15 : rom_data_pri =  150'b000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000;
		8'd16 : rom_data_pri =  150'b000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000;
		8'd17 : rom_data_pri =  150'b000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000;
		8'd18 : rom_data_pri =  150'b000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000;
		8'd19 : rom_data_pri =  150'b000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000;
		8'd20 : rom_data_pri =  150'b000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000;
		8'd21 : rom_data_pri =  150'b000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000;
		8'd22 : rom_data_pri =  150'b000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
		8'd23 : rom_data_pri =  150'b000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000;
		8'd24 : rom_data_pri =  150'b000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000;
		8'd25 : rom_data_pri =  150'b000000000000110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001000000000000;
		8'd26 : rom_data_pri =  150'b000000000000111001111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111000011000000000000;
		8'd27 : rom_data_pri =  150'b000000000000111100111100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000111000000000000;
		8'd28 : rom_data_pri =  150'b000000000000011110001111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011110001110000000000000;
		8'd29 : rom_data_pri =  150'b000000000000011111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111100111110000000000000;
		8'd30 : rom_data_pri =  150'b000000000000001100110011110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001111001111100000000000000;
		8'd31 : rom_data_pri =  150'b000000000000000110011001111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011100011001100000000000000;
		8'd32 : rom_data_pri =  150'b000000000000000011001100111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100111000100111000000000000000;
		8'd33 : rom_data_pri =  150'b000000000000000011100100001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110011001110000000000000000;
		8'd34 : rom_data_pri =  150'b000000000000000000010000000010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001000000011000000000000000000;
		8'd35 : rom_data_pri =  150'b000000000000000000011011110000011100000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011100110000000000000000000;
		8'd36 : rom_data_pri =  150'b000000000000000111001011111100001110000000000000000000000000000000000000000000111000000000000000000000000000000000011100000111110100011000000000000000;
		8'd37 : rom_data_pri =  150'b000000000000000111100001111111001111100000000000000000000000000000000000001111111100000000000000000000000000000000111100011111110001111000000000000000;
		8'd38 : rom_data_pri =  150'b000000000000000011110000110011100111110000000000000000000000000000000000011111111100000000000000000000000000000011111001111011100011111000000000000000;
		8'd39 : rom_data_pri =  150'b000000000000000011111100011001110011111000000000000000000000000000000000111111111110000000000000000000000000000111110011110111000111110000000000000000;
		8'd40 : rom_data_pri =  150'b000000000000000001111111001100011000111110000000000000000000000000000001111111111110000000000000000000000000001111100111001110011111110000000000000000;
		8'd41 : rom_data_pri =  150'b000000000000000000111111000110001100111111100000000000000000000000000000111111111111000000000000000000000000111111001110011000111111100000000000000000;
		8'd42 : rom_data_pri =  150'b000000000000000000011111110011100110001111110000000000000000000000000001111111111111000000000000000000000001111110011000110001111111000000000000000000;
		8'd43 : rom_data_pri =  150'b000000000000000000000101111000110000000111111100000000000000000000000001111111111111000000000000000000000111111000010011100111111100000000000000000000;
		8'd44 : rom_data_pri =  150'b000000000000000000000110111100001100110011111110000000000000000000000001111111111111100000000000000000001111110001000110001111011000000000000000000000;
		8'd45 : rom_data_pri =  150'b000000000000000000000111001111000100111100111111000000000000000000000001111111111111100000000000000000111111100111001100011110011000000000000000000000;
		8'd46 : rom_data_pri =  150'b000000000000000000000011100111100000111111111111110000000000000000000011111111111111100000000000000001111110011111000001111000110000000000000000000000;
		8'd47 : rom_data_pri =  150'b000000000000000000000001110011101100011111111111111000000000000000000011111111111111100000000000000011111111111110000101110001100000000000000000000000;
		8'd48 : rom_data_pri =  150'b000000000000000000000000111100111110000111111111111100000000000000000011111111111111100000000000000111111111111100011111100111000000000000000000000000;
		8'd49 : rom_data_pri =  150'b000000000000000000000000011110001111000011111111111110000000000000000011111111111111110000000000001111111111111000111110001110000000000000000000000000;
		8'd50 : rom_data_pri =  150'b000000000000000000000000000111000011011001111111111110000000000000000011111111111111100000000000011111111111100000111000111100000000000000000000000000;
		8'd51 : rom_data_pri =  150'b000000000000000000000010000011110000011100111111111111000000000000000111111111111111110000000000111111111111001110000011110000000000000000000000000000;
		8'd52 : rom_data_pri =  150'b000000000000000000000011111000111110001111111111111111000000000000000111111111111111110000000000111111111111111100001111100001111000000000000000000000;
		8'd53 : rom_data_pri =  150'b000000000000000000000011111100000001100111111111111111000000000000000111111111111111100000000000111111111111111000111100001111110000000000000000000000;
		8'd54 : rom_data_pri =  150'b000000000000000000000000011110100001110011111111111111100000000000000111111111111111100000000000111111111111110001100000011110000000000000000000000000;
		8'd55 : rom_data_pri =  150'b000000000000000000000000011100111000011001111111111111000000000000000111111111111111100000000000111111111111100111000011001110000000000000000000000000;
		8'd56 : rom_data_pri =  150'b000000000000000000000000010110111110000000011111111111000000000000001111111111111111110000000000111111111111000000001111001111000000000000000000000000;
		8'd57 : rom_data_pri =  150'b000000000000000000000000000010011111100111111111111111000000000000001111111111111111110000000000111111111110011001111110010000000000000000000000000000;
		8'd58 : rom_data_pri =  150'b000000000000000000000000000111001000110011111111111111000000000000001111111111111111110000000000011111111111110011110010011000000000000000000000000000;
		8'd59 : rom_data_pri =  150'b000000000000000000000000000011100110000001111111111110000000000000001111111111111111110000000000011111111111100100000100110000000000000000000000000000;
		8'd60 : rom_data_pri =  150'b000000000000000000000000000001110001100000011111111100000000000000001111111111111111110000000000001111111111000000110001100000000000000000000000000000;
		8'd61 : rom_data_pri =  150'b000000000000000000000000000000011000011111000111111110000000000001111111111111111111110000000000001111111100011111000011000000000000000000000000000000;
		8'd62 : rom_data_pri =  150'b000000000000000000000000000000000111000000000001111110000000000011111111111111111111110000000000011111100000100000011100000000000000000000000000000000;
		8'd63 : rom_data_pri =  150'b000000000000000000000000000000110000111110011111111111000000000011111111111111111111110000000000011111100110000011100001000000000000000000000000000000;
		8'd64 : rom_data_pri =  150'b000000000000000000000000000000011100000000001111111111111100000111111111111111111111110000000000111111111100111000000111000000000000000000000000000000;
		8'd65 : rom_data_pri =  150'b000000000000000000000000000000011111110000100001000111111111100111111111111111111111111001111111111111111000000000111110000000000000000000000000000000;
		8'd66 : rom_data_pri =  150'b000000000000000000000000000000001111100111100000001111111111100111111111111111111111111100111111111100000011110011111100000000000000000000000000000000;
		8'd67 : rom_data_pri =  150'b000000000000000000000000000000000111100110001110011111111111100111111111111111111111111100111111111111010000011001111000000000000000000000000000000000;
		8'd68 : rom_data_pri =  150'b000000000000000000000000000000000001100000000000000111101111100111111111111111111111111100111111111100000111011001110000000000000000000000000000000000;
		8'd69 : rom_data_pri =  150'b000000000000000000000000000000000000111000000001100000001111100111111111111111111111111100111100000001100000000011000000000000000000000000000000000000;
		8'd70 : rom_data_pri =  150'b000000000000000000000000000000000000001111111011110000111111100111111111111111111111111100111111000011100111111110000000000000000000000000000000000000;
		8'd71 : rom_data_pri =  150'b000000000000000000000000000000000000000000100010000110001100100111111111111111111111111110011110011000110011110000000000000000000000000000000000000000;
		8'd72 : rom_data_pri =  150'b000000000000000000000000000000000000000000000011111000100000000111111111111111111111111110000000001110111000000000000000000000000000000000000000000000;
		8'd73 : rom_data_pri =  150'b000000000000000000000000000000000000001111111000000000110110000111111111111111111111111110010001000000000000001100000000000000000000000000000000000000;
		8'd74 : rom_data_pri =  150'b000000000000000000000000000000000000001111100000111110110110000111111111111111111111111100011111011000000111111100000000000000000000000000000000000000;
		8'd75 : rom_data_pri =  150'b000000000000000000000000000000000000000110000011111000011111100111111111111111111111111100011111001111100000011100000000000000000000000000000000000000;
		8'd76 : rom_data_pri =  150'b000000000000000000000000000000000000000011111111100001000011000111111111111111111111111100110000000011111110111000000000000000000000000000000000000000;
		8'd77 : rom_data_pri =  150'b000000000000000000000000000000000000000000110000000010000000000111111111111111111111111100110000110000011111100000000000000000000000000000000000000000;
		8'd78 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000111010100000100111111111111111111111111100000011010110000000000000000000000000000000000000000000000000;
		8'd79 : rom_data_pri =  150'b000000000000000000000000000000000000000000000111111011001001110111111111111111111111111100100101010111110000000000000000000000000000000000000000000000;
		8'd80 : rom_data_pri =  150'b000000000000000000000000000000000000000000000011111010011001100011111111111111111111111100100110110111111000000000000000000000000000000000000000000000;
		8'd81 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000111100000011111111111111111111111100101111000111100000000000000000000000000000000000000000000000;
		8'd82 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111111011100001110000000000000000000000000000000000000000000000000000000;
		8'd83 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111110011110000000000000000000000000000000000000000000000000000000000000;
		8'd84 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111110011110000000000000000000000000000000000000000000000000000000000000;
		8'd85 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111110011110000000000000000000000000000000000000000000000000000000000000;
		8'd86 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011100111111111111110011110000000000000000000000000000000000000000000000000000000000000;
		8'd87 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111110011110000000000000000000000000000000000000000000000000000000000000;
		8'd88 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111110001110000000000000000000000000000000000000000000000000000000000000;
		8'd89 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111111001111000000000000000000000000000000000000000000000000000000000000;
		8'd90 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111111001111000000000000000000000000000000000000000000000000000000000000;
		8'd91 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111111111111000000000000000000000000000000000000000000000000000000000000;
		8'd92 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111111111111000000000000000000000000000000000000000000000000000000000000;
		8'd93 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'd94 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111100111111111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'd95 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111000111111111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'd96 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111100000000000000000000000000000000000000000000000000000000000;
		8'd97 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111110000000000000000000000000000000000000000000000000000000000;
		8'd98 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111110000000000000000000000000000000000000000000000000000000000;
		8'd99 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111110000000000000000000000000000000000000000000000000000000000;
		8'd100 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111110000000000000000000000000000000000000000000000000000000000;
		8'd101 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111111000000000000000000000000000000000000000000000000000000000;
		8'd102 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111111000000000000000000000000000000000000000000000000000000000;
		8'd103 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111111000000000000000000000000000000000000000000000000000000000;
		8'd104 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111111100000000000000000000000000000000000000000000000000000000;
		8'd105 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111001111111111111111111111111100000000000000000000000000000000000000000000000000000000;
		8'd106 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000110011111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'd107 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'd108 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'd109 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'd110 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'd111 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'd112 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000;
		8'd113 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111111111111111000111111111111110000000000000000000000000000000000000000000000000000000;
		8'd114 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111111111111110000011111111111110000000000000000000000000000000000000000000000000000000;
		8'd115 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111111111111100000001111111111110000000000000000000000000000000000000000000000000000000;
		8'd116 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111111111111000000001111111111110000000000000000000000000000000000000000000000000000000;
		8'd117 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000000111111111110000000001111111111110000000000000000000000000000000000000000000000000000000;
		8'd118 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000001111111111110000000000111111111110000000000000000000000000000000000000000000000000000000;
		8'd119 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000001111111111100000000000111111111110000000000000000000000000000000000000000000000000000000;
		8'd120 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000001111111111100000000000011111111110000000000000000000000000000000000000000000000000000000;
		8'd121 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000001111111111000000000000011111111110000000000000000000000000000000000000000000000000000000;
		8'd122 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000001111111110000000000000001111111110000000000000000000000000000000000000000000000000000000;
		8'd123 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000001111111110000000000000000111111110000000000000000000000000000000000000000000000000000000;
		8'd124 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000;
		8'd125 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111000000000000000000000000000000000000000000000000000000;
		8'd126 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000;
		8'd127 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000;
		8'd128 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000;
		8'd129 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111100000000000000000000000000000000000000000000000000000;
		8'd130 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000001111111110000000000000000000001111111110000000000000000000000000000000000000000000000000000;
		8'd131 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000111111110000000000000000000000000000000000000000000000000000;
		8'd132 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000111111110000000000000000000000000000000000000000000000000000;
		8'd133 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000011111110000000000000000000000000000000000000000000000000000;
		8'd134 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000011111111000000000000000000000000000000000000000000000000000;
		8'd135 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000011111111000000000000000000000000000000000000000000000000000;
		8'd136 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000001111111100000000000000000000000000000000000000000000000000;
		8'd137 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000001111111100000000000000000000000000000000000000000000000000;
		8'd138 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000111111110000000000000000000000000000000000000000000000000;
		8'd139 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000;
		8'd140 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000011111111000000000000000000000000000000000000000000000000;
		8'd141 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000011111111000000000000000000000000000000000000000000000000;
		8'd142 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001111111000000000000000000000000000000000000000000000000;
		8'd143 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000001111111100000000000000000000000000000000000000000000000;
		8'd144 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000111111100000000000000000000000000000000000000000000000;
		8'd145 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000;
		8'd146 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000;
		8'd147 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000;
		8'd148 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000;
		8'd149 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000;
		8'd150 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000;
		8'd151 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000;
		8'd152 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000;
		8'd153 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000;
		8'd154 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000;
		8'd155 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000;
		8'd156 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000;
		8'd157 : rom_data_pri =  150'b000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000;
		8'd158 : rom_data_pri =  150'b000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000;
		8'd159 : rom_data_pri =  150'b000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000;
		8'd160 : rom_data_pri =  150'b000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000;
		8'd161 : rom_data_pri =  150'b000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000;
		8'd162 : rom_data_pri =  150'b000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000;
		8'd163 : rom_data_pri =  150'b000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000;
		8'd164 : rom_data_pri =  150'b000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000;
		8'd165 : rom_data_pri =  150'b000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000;
		8'd166 : rom_data_pri =  150'b000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000;
		8'd167 : rom_data_pri =  150'b000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000;
		8'd168 : rom_data_pri =  150'b000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000;
		8'd169 : rom_data_pri =  150'b000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000;
		8'd170 : rom_data_pri =  150'b000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000;
		8'd171 : rom_data_pri =  150'b000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000;
		8'd172 : rom_data_pri =  150'b000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000;
		8'd173 : rom_data_pri =  150'b000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000;
		8'd174 : rom_data_pri =  150'b000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000;
		8'd175 : rom_data_pri =  150'b000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000;
		8'd176 : rom_data_pri =  150'b000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001100100000000000000000000000000000000000000;
		8'd177 : rom_data_pri =  150'b000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
		8'd178 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001000110000000000000000000000000000000000000;
		8'd179 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001110110000000000000000000000000000000000000;
		8'd180 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000;
		8'd181 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000;
		8'd182 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000;
		8'd183 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000;
		8'd184 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000;
		8'd185 : rom_data_pri =  150'b000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000;
		8'd186 : rom_data_pri =  150'b000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

	endcase
	
	//-----------------------------PRINCESS-----------------------------			
			
	assign pri_x_l = pri_x_reg;
	assign pri_y_t = 230;
	assign pri_x_r  = pri_x_l  + PRI_LO_SIZE - 1;
	assign pri_y_b  = pri_y_t  + PRI_HI_SIZE - 1; 
	assign sq_pri_on =pri_turn_reg&& (pri_x_l <= pix_x) && (pix_x <= pri_x_r) && (pri_y_t <= pix_y)  && (pix_y <= pri_y_b);
	//draw detail of princess
	assign rom_addr_pri  = pix_y [7:0] - pri_y_t[7:0] ; 
	assign rom_col_pri  = pix_x [7:0] - pri_x_l[7:0] ; 
	assign rom_bit_pri  = rom_data_pri [rom_col_pri] ; 
	assign rd_pri_on  = sq_pri_on & rom_bit_pri;
	
	//update position for princess
	always@*			
		begin				
			begin
				pri_x_next = pri_x_reg;					
				if(pri_turn_reg&refr_tick & ~KEY[0] & at_mid_reg )
					pri_x_next = pri_x_reg - mario_del_run_next;
				end
		end

//-------------------------------------------------MOUNTAIN----------------------------------------------------------
	localparam mtn_LO_SIZE = 273;
	localparam mtn_HI_SIZE = 94;
	reg [9:0] mtn_x_reg;
	reg [9:0] mtn_x_next;
	wire [9:0]mtn_x_l,mtn_x_r;
	wire [9:0]mtn_y_t,mtn_y_b; 
		//draw mountain
	wire [6:0] rom_addr_mtn;
	wire [8:0] rom_col_mtn;
	reg [273:0] rom_data_mtn;
	wire rom_bit_mtn;
	wire sq_mtn_on, rd_mtn_on;
	reg [8:0] mtn_rgb = 9'b111111111;
	
	always @*
	case(rom_addr_mtn)

		7'd0: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd1: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd2: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd3: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd4: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd5: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd6: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd7: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd8: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd9: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd10: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd11: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd12: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd13: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd14: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd15: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd16: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd17: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000001111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd18: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000001111100000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd19: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000111111000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd20: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000011111000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000;
		7'd21: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000111111000000000000000111110000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000001111111111111111110010000000000000000000000000000000000000000000000000000000000000000000;
		7'd22: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000011111110000000000000000011111000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000;
		7'd23: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000111111100000000000000000011111110000000000000000000100000000000000011111111111111111100000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000;
		7'd24: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000001111110000000000000000000000011111000000000000000001100000000000000111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111110000000000011000000000000000000000000000000000000000000000000;
		7'd25: rom_data_mtn = 274'b000000000000000000000000000000000111000000000000000111111000000000000000000000000011111110000000000001111110000000000011111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111100000000000111100000000000000000000000000000000000000000000000;
		7'd26: rom_data_mtn = 274'b000000000000000000000000000000000011100000000000001111110000000000000000000000000000111110000000000111111110000000011111111111111111111111111111100000000000000000000000000000000000001111111111111111111111111111000000000011111110000000000000000000000000000000000000000000000;
		7'd27: rom_data_mtn = 274'b000000000000000000000000000000000101111000000000011111000000000000000000000000000000011111000000111111111111110000111111111111111111111111111111111000000000000000000000000000000000001111111111111111111111110000000000000111111111110000000000000000000000000000000000000000000;
		7'd28: rom_data_mtn = 274'b000000000000000000000000000000011100011110000001111111000000000000000000000000000000000111110111111111100001111111111111111111111111111111111111111111111000000000000000000000000000000001111001111111111111000000000000011111000111110000000000000000000000000000000000000000000;
		7'd29: rom_data_mtn = 274'b000000000000000000000000000000111100000111111111111000000000000000000000000000000000000001111111111100000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111100000011111100000000000000000000000000000000000000000;
		7'd30: rom_data_mtn = 274'b000000000000000000000000000001111100000001111111110000000000000000000000000000000000000000111111100000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111100000000011110000000000000000000000000000000000000000;
		7'd31: rom_data_mtn = 274'b000000000000000000000000000001100000000000011111100000000000000000000000000000000000000000011111000000011111111111111111101111111111111111111110001111111111100000000000000000000000000000000000000000000000000000000111111000000000011111000000000000000000000000000000000000000;
		7'd32: rom_data_mtn = 274'b000000000000000000000000000011100000000000001111000000000000000000000000000000000000000000011110000011111111111110000100000001111111111111110000000011111111111000000000000000000000000000000000000000000000000000001111100000000000001111100000000000000000000000000000000000000;
		7'd33: rom_data_mtn = 274'b000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000011111111111100000000000001111111110000000000000000000000000000000000000000000000000011111000000000000000011111000000000000000000000000000000000000;
		7'd34: rom_data_mtn = 274'b000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000111111000000000000000000111111111100000000000000000000000000000001000000000001110111110000000000000000011111100000000000000000000000000000000000;
		7'd35: rom_data_mtn = 274'b000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000001110000000000000000000001111111111111000000000000000000000000001100000011111111111000000000000000000001111110000000000000000000000000000000000;
		7'd36: rom_data_mtn = 274'b000000000000000000000111110000000000000000000000001111000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000001111111111100000000000000000000001111110000111111111110000000000000000000000001111000000000000111000000000000000000;
		7'd37: rom_data_mtn = 274'b000000000000000000001111100000000000000000000000011111110000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000001111011111111111111111000000000000000000000000111111000000001111000000000000000000;
		7'd38: rom_data_mtn = 274'b000000000000000011111110000000000000000000000000111111111110000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000001001111111111111111111110000000000000000000000011111100001111001111000000000000000;
		7'd39: rom_data_mtn = 274'b000000000000000111111100000000000000000000000001111111111111110000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000111111111111111111111111111100000000000000000000001111101111110001111000000000000000;
		7'd40: rom_data_mtn = 274'b000000000000001111111000000000000000000000001111111111111111111100000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111111111111111111111111111111000000000000000000000111111110000000001100000000000000;
		7'd41: rom_data_mtn = 274'b000000000000001111110000000000000000000000011111111111111111111111111110000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110111111111111111111111111000000000000000000000111000000000001100000000000000;
		7'd42: rom_data_mtn = 274'b000000000000000100000000000000000000000001111111111111111111100011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111000000011110000000110011111100000000000000000000000000000000000111000000000000;
		7'd43: rom_data_mtn = 274'b000000000000000000000000000000000000000111111110000111111110000000001111111111111111100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000011111100000000000000000000000000000000011110000000000;
		7'd44: rom_data_mtn = 274'b000000000000000000000000000000000000011111100000000000001000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000011111100000000000000000000000000000011111000000000;
		7'd45: rom_data_mtn = 274'b000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000111110000000000000000000000000000000111110000000;
		7'd46: rom_data_mtn = 274'b000000000000000000000000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000001111110000;
		7'd47: rom_data_mtn = 274'b000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000111111000;
		7'd48: rom_data_mtn = 274'b000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000011111111;
		7'd49: rom_data_mtn = 274'b000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000011100;
		7'd50: rom_data_mtn = 274'b000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000;
		7'd51: rom_data_mtn = 274'b000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000;
		7'd52: rom_data_mtn = 274'b000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000;
		7'd53: rom_data_mtn = 274'b000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000;
		7'd54: rom_data_mtn = 274'b000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000;
		7'd55: rom_data_mtn = 274'b000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000;
		7'd56: rom_data_mtn = 274'b000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd57: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd58: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd59: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000;
		7'd60: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000;
		7'd61: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000;
		7'd62: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000;
		7'd63: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000111100000000000000000000000000000000000000000000;
		7'd64: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000111100000000000000000000000000000000000000000000;
		7'd65: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111100000111100000000000000000000000000000000000000000000;
		7'd66: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111100000111100000000000000000000000000000000000000000000;
		7'd67: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110011111111100001111110000000000000000000000000000000000000000000;
		7'd68: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110011111111100001111110000000000000000000000000000000000000000000;
		7'd69: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011111111111011111110000000000000000000000000000000000000000000;
		7'd70: rom_data_mtn = 274'b000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011111111111011111110000000000000000000000000000000000000000000;
		7'd71: rom_data_mtn = 274'b000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000110000011111110000000000000000000000000000000000000000000;
		7'd72: rom_data_mtn = 274'b000000000000000000000000000000000000000010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100010001000111110000000110000000110000000000000000000000000000000000000000000000;
		7'd73: rom_data_mtn = 274'b000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000110000100000000000000000000000000000000000000000000000000000000;
		7'd74: rom_data_mtn = 274'b000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111100000001010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000;
		7'd75: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010100000000000000000000000;
		7'd76: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000110000000000000000000;
		7'd77: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111111111111111111111111110000000000000000000;
		7'd78: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd79: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000;
		7'd80: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd81: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111111111111111111111111111111111111111000000000000000000;
		7'd82: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000000000;
		7'd83: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd84: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd85: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd86: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd87: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd88: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd89: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd90: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd91: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd92: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd93: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		7'd94: rom_data_mtn = 274'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	endcase

	//-----------------------------MOUNTAIN 1-----------------------------			
		
	assign mtn_x_l = mtn_x_reg;
	assign mtn_y_t = 336;
	assign mtn_x_r  = mtn_x_l  + mtn_LO_SIZE - 1;
	assign mtn_y_b  = mtn_y_t  + mtn_HI_SIZE - 1; 
	assign sq_mtn_on = (mtn_x_l <= pix_x) && (pix_x <= mtn_x_r) && (mtn_y_t <= pix_y)  && (pix_y <= mtn_y_b);
	//draw detail of mountain
	assign rom_addr_mtn  = pix_y [6:0] - mtn_y_t[6:0] ; //3bits
	assign rom_col_mtn  = pix_x [8:0] - mtn_x_l[8:0] ; //1 bit
	assign rom_bit_mtn  = rom_data_mtn [rom_col_mtn] ; 
	assign rd_mtn_on  = sq_mtn_on & rom_bit_mtn;
	
	//update position of mountain
	always@*			
		begin
			mtn_x_next = mtn_x_reg;
			if(refr_tick & ~KEY[0] & at_mid_reg )
				mtn_x_next = mtn_x_reg - mario_del_run_next;
		end		
	
	
	//--------------------------WALL--------------------------------
	
	localparam wall_hi_size = 32;
	reg [9:0]wall_lo_size_reg ;
	reg [9:0]wall_lo_size_next;
	wire [9:0] wall_x_l, wall_x_r, wall_y_b, wall_y_t;
	reg [9:0]wall_x_next;	
	reg [9:0]wall_x_reg;
	reg [9:0]wall_y_next;	
	reg [9:0]wall_y_reg;
	wire wall_black;
	assign wall_black = wall_x_l<=pix_x && pix_x<=wall_x_r && pix_y<=wall_y_b && pix_y>=wall_y_t; //the background of wall
	wire wall_on;
	reg [8:0]wall_rgb = 9'b011001000; //black

	
	//--------------------------CLOULD---------1-----------------------------------
	localparam C1_LO_SIZE = 116;
	localparam C1_HI_SIZE = 39;
	reg [9:0] c1_x_reg;
	reg [9:0] c1_x_next;
	wire [9:0] c1_x_l, c1_x_r;
	wire [9:0] c1_y_t, c1_y_b; 
	//--------------------------DRAW CLOULD--------1-----------------------------------
	wire [5:0] rom_addr_c1;
	wire [6:0] rom_col_c1;
	reg [115:0] rom_data_c1;
	wire rom_bit_c1;
	wire sq_c1_on, rd_c1_on;
	reg [8:0] c1_rgb = 9'b111111111;
	
	always @*
	case(rom_addr_c1)
	
			6'd0: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000;
			6'd1: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000;
			6'd2: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000;
			6'd3: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000;
			6'd4: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000;
			6'd5: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000;
			6'd6: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000111111100000000000000000;
			6'd7: rom_data_c1 = 116'b  00000000000000000000000000000000000000000000000000000000001111111111111111111111111111110011111111111000000000000000;
			6'd8: rom_data_c1 = 116'b  00000000000000000000000000000000000000000111111100000000001111111111111111111111111111111111111111111110000000000000;
			6'd9: rom_data_c1 = 116'b  00000000000000000000000000000000000001111111111111111000000011111111111111111111111111111111111111111111000000000000;
			6'd10: rom_data_c1 = 116'b 00000000000000000000000000000000001111111111111111111111000000111111111111111111111111111111111111111111100000000000;
			6'd11: rom_data_c1 = 116'b 00000000000000000000000000000000111111111111111111111111110000001111111111111111111111111111111111111111100000000000;
			6'd12: rom_data_c1 = 116'b 00000000000000000000000000000011111111111111111111111111111100000111111111111111111111111111111111111111100000000000;
			6'd13: rom_data_c1 = 116'b 00000000000000000000000000001111111111111111111111111111111111000001111111111111111111111111111111111111111111111110;
			6'd14: rom_data_c1 = 116'b 00000000000000000000000000011111111111111111111111111111111111100000111111111111111111111111111111111111111111111111;
			6'd15: rom_data_c1 = 116'b 00000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000;
			6'd16: rom_data_c1 = 116'b 00000000000000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000;
			6'd17: rom_data_c1 = 116'b 00000000000000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000;
			6'd18: rom_data_c1 = 116'b 00000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000;
			6'd19: rom_data_c1 = 116'b 00000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000;
			6'd20: rom_data_c1 = 116'b 00000000000000000000001111111111111111111111111111111111111111111110000000011111111111111000000000000000000000000000;
			6'd21: rom_data_c1 = 116'b 00000000000000000000001111111111111111111111111111111111111111111111000111111111111111111111000000000000000000000000;
			6'd22: rom_data_c1 = 116'b 00000000000000000000001111111111111111111111111111111111111111111111001111111111111111111111110000000000000000000000;
			6'd23: rom_data_c1 = 116'b 00000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000;
			6'd24: rom_data_c1 = 116'b 00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000;
			6'd25: rom_data_c1 = 116'b 00000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000;
			6'd26: rom_data_c1 = 116'b 00000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000;
			6'd27: rom_data_c1 = 116'b 00000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
			6'd28: rom_data_c1 = 116'b 00000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
			6'd29: rom_data_c1 = 116'b 00000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
			6'd30: rom_data_c1 = 116'b 00000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
			6'd31: rom_data_c1 = 116'b 00000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
			6'd32: rom_data_c1 = 116'b 00001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000;
			6'd33: rom_data_c1 = 116'b 00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000;
			6'd34: rom_data_c1 = 116'b 00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000;
			6'd35: rom_data_c1 = 116'b 01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100;
			6'd36: rom_data_c1 = 116'b 11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
			6'd37: rom_data_c1 = 116'b 11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			6'd38: rom_data_c1 = 116'b 00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
		
	endcase
	
	//-----------------------------CLOUD_ 1-----------------------------			
			
	assign c1_x_l = c1_x_reg;
	assign c1_y_t = 150;
	assign c1_x_r  = c1_x_l  + C1_LO_SIZE - 1;
	assign c1_y_b  = c1_y_t  + C1_HI_SIZE - 1; 
	assign sq_c1_on = (c1_x_l <= pix_x) && (pix_x <= c1_x_r) && (c1_y_t <= pix_y)  && (pix_y <= c1_y_b);
	
	assign rom_addr_c1  = pix_y [5:0] - c1_y_t[5:0] ; //3bits
	assign rom_col_c1  = pix_x [6:0] - c1_x_l[6:0] ; //1 bit
	assign rom_bit_c1  = rom_data_c1 [rom_col_c1] ; 
	assign rd_c1_on  = sq_c1_on & rom_bit_c1;
	
	//update the position of cloud
	always@*			
		begin
			c1_x_next = c1_x_reg;
			if(refr_tick & ~KEY[0] & at_mid_reg )
				c1_x_next = c1_x_reg - mario_del_run_next;
		end		
		
	
	//--------------------------CLOULD-----------------------------------
	localparam C_LO_SIZE = 64;
	localparam C_HI_SIZE = 16;
	reg [9:0] c_x_reg;
	reg [9:0] c_x_next;
	wire [9:0] c_x_l, c_x_r;
	wire [9:0] c_y_t, c_y_b; 
	//draw detail of cloud
	wire [3:0] rom_addr_c;
	wire [5:0] rom_col_c;
	reg [63:0] rom_data_c;
	wire rom_bit_c;
	wire sq_c_on, rd_c_on;
	reg [8:0] c_rgb = 9'b111111111;
	
	//-------------------------- DRAW WALLL-----------------------------------
	wire [4:0] rom_addr_w;
	wire [7:0] rom_col_w;
	reg [299:0] rom_data_w;
	wire rom_bit_w;
	wire rd_wall_on;

	always @*
	case(rom_addr_c)
	
		4'd0 : rom_data_c =  64'b0000000000000000000000000000001111111111100000000000000000000000;                      
		4'd1 : rom_data_c =  64'b0000000000000000000000001111111111111111111110000000000000000000;                  
		4'd2 : rom_data_c =  64'b0000000000000000000000111111111111111111111111100000000000000000;                
		4'd3 : rom_data_c =  64'b0000000000000000000011111111111111111111111111110000000000000000;               
		4'd4 : rom_data_c =  64'b0000000000000011111111111111111111111111111111111000000000000000;             
		4'd5 : rom_data_c =  64'b0000000000000111111111111111111111111111111111111100000000000000;             
		4'd6 : rom_data_c =  64'b0000001111111111111111111111111111111111111111111111110000000000;         
		4'd7 : rom_data_c =  64'b0011111111111111111111111111111111111111111111111111111111111000;  
		4'd8 : rom_data_c =  64'b0111111111111111111111111111111111111111111111111111111111111110;
		4'd9 : rom_data_c =  64'b0111111111111111111111111111111111111111111111111111111111111110;
		4'd10: rom_data_c =  64'b1111111111111111111111111111111111111111111111111111111111111111;
		4'd11: rom_data_c =  64'b0111111111111111111111111111111111111111111111111111111111111111;
		4'd12: rom_data_c =  64'b0111111111111111111111111111111111111111111111111111111111111110;
		4'd13: rom_data_c =  64'b0001111111111111111111111111111111111111111111111111111111111100; 
		4'd14: rom_data_c =  64'b0000000111111111111111111111111111111111111111111111111111000000;       
		4'd15: rom_data_c =  64'b0000000000000111111111111111111111111111111111111111111000000000;
	endcase


	//Rom memory for drawing detail of brick (wall)
	always@*
	case(rom_addr_w)
		5'd0 : rom_data_w =  300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd1 : rom_data_w =  300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd2 : rom_data_w =  300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd3 : rom_data_w =  300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd4 : rom_data_w =  300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd5 : rom_data_w =  300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd6 : rom_data_w =  300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd7 : rom_data_w =  300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd8 : rom_data_w =  300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd9 : rom_data_w =  300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd10 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd11 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd12 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd13 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd14 : rom_data_w = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd15 : rom_data_w = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd16 : rom_data_w = 300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd17 : rom_data_w = 300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd18 : rom_data_w = 300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd19 : rom_data_w = 300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd20 : rom_data_w = 300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd21 : rom_data_w=  300'b111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111001;
		5'd22 : rom_data_w = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd23 : rom_data_w = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd24 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd25 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd26 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd27 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd28 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd29 : rom_data_w = 300'b111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111111111110001111111111111111111111000111111111111111111111100011111111111111;
		5'd30 : rom_data_w = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		5'd31 : rom_data_w = 300'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;		
		 
	endcase
	
	
	//-----------------------------------PIPE1------------------------------------
	
	localparam pipe1_lo_size = 71; //pipe1 long size
	localparam pipe1_hi_size = 64; //pipe1 high size
	localparam pipe1_y_t = BASE - pipe1_hi_size; //base always stand on Ground	
	wire [9:0] pipe1_x_l, pipe1_x_r, pipe1_y_b;
	reg [9:0] pipe1_x_reg, pipe1_x_next;
	wire pipe1_on;
	reg [8:0]pipe1_rgb = 9'b000011000; //Green color	
	//draw pipe
	wire [5:0] rom_addr_p1;
	wire [6:0] rom_col_p1;
	reg [70:0] rom_data_p1;
	wire rom_bit_p1;
	wire rd_p1_on;
		
	always@*
		case(rom_addr_p1)

		6'd0 :rom_data_p1  =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd3 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd4 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd5 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd6 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd7 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd8 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd9 : rom_data_p1 =  71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd10 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd11 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd12 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd13 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
	    6'd14 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
	    6'd15 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
	    6'd16 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
	    6'd17 : rom_data_p1 = 71'b11111111111111111111111111111111111111111111111111111111111111111111111;
		6'd18 : rom_data_p1 = 71'b00000111000000000000000000000000000000000000000000000000000000011100000;
		6'd19 : rom_data_p1 = 71'b00000111000000000000000000000000000000000000000000000000000000011100000;
	    6'd20 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;   
        6'd21 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
	    6'd22 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd23 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd24 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd25 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd26 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd27 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd28 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd29 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd30 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd31 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd32 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd33 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd34 : rom_data_p1 = 71'b00000111111111111111111111111111111111111111110100111111111111111100000;
		6'd35 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd36 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd37 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd38 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd39 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd40 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd41 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd42 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd43 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd44 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd45 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd46 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd47 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd48 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd49 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd50 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd51 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd52 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd53 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd54 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd55 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd56 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd57 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd58 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd59 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
		6'd60 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;											   
        6'd61 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000 ;   
		6'd62 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
        6'd63 : rom_data_p1 = 71'b00000111111111111111111111111111111111110011110100111111111111111100000;
	endcase
	
		//Reading pixel in rom memory
	    assign rom_addr_p1  = pix_y [5:0] - pipe1_y_t[5:0] ; //3bits
		assign rom_col_p1  = pix_x [6:0] - pipe1_x_l[6:0] ; //1 bit
		assign rom_bit_p1  = rom_data_p1 [rom_col_p1] ; 
		assign rd_p1_on  = rd_pipe1_on & rom_bit_p1;	
	
	//-----------------------------------HOLE------------------------------------
	
	localparam hole1_lo_size = 100;	
	localparam hole1_hi_size = 50 + 1;	
	
	wire [9:0] hole1_x_l, hole1_x_r, hole1_y_b, hole1_y_t;
	reg [9:0] hole1_x_reg, hole1_x_next;
	wire hole1_on;
	wire [8:0] hole1_rgb;
	//--------------------------------------------monster(DRAGON)----------------------------------------------
	localparam MONSTER_X = 76;
	localparam MONSTER_Y = 71;
	reg mst_turn_reg;
    reg mst_turn_next;
	wire [9:0] monster_x_l, monster_x_r, monster_y_t, monster_y_b;
	reg [9:0] monster_x_reg, monster_y_reg;
	wire [9:0] monster_x_next, monster_y_next;
	reg  [9:0]  mstX_delta_reg , mstX_delta_next ; 
	reg  [9:0]  mstY_delta_reg,  mstY_delta_next;
	localparam  MONSTER_V_P = 2;
	localparam  MONSTER_V_N = -2; 
	wire monster_on;
	wire [8:0] monster_rgb; 
	//--------------------------MUSHROOM--------------------------------

	localparam mushroom_lo_size = 25;
	localparam mushroom_hi_size = 25;
	
	wire [9:0]mushroom_x_next,mushroom_y_next;
	reg [9:0]mushroom_x_reg,mushroom_y_reg;	
	wire [9:0] mushroom_x_l,mushroom_x_r,mushroom_y_t,mushroom_y_b;	
	
	wire sq_mushroom_on;
	reg [9:0] mushroom_rgb = 9'b111101000;//RED
	wire [2:0] mushroom_stage_next;
	reg	[2:0] mushroom_stage_reg; //stage = 1: right | 2: left | 3: up | 4: down |5: back to base | 6: begin | 7 : disappear
	assign mushroom_x_l = mushroom_x_reg;
	assign mushroom_y_t = mushroom_y_reg;	
	assign mushroom_x_r = mushroom_x_l + mushroom_lo_size;
	assign mushroom_y_b = mushroom_y_t + mushroom_hi_size;		
	assign sq_mushroom_on = ( mushroom_x_l <= pix_x ) && (pix_x <= mushroom_x_r) && (mushroom_y_t <= pix_y) && (pix_y <= mushroom_y_b);
	//moving of mushroom
	assign mushroom_x_next 	= (refr_tick && mushroom_stage_reg==6) ?(wall_x_l+25) // 6: begin
				: (refr_tick &&  mushroom_stage_reg==7) ? 639					// 7 : disappear
				: (refr_tick && mushroom_stage_reg==1) ? (mushroom_x_reg + 1) 			//1: right
				: (refr_tick && mushroom_stage_reg==2) ? (mushroom_x_reg - 1)	 		//  2:left
				: (mushroom_x_reg);
	assign mushroom_y_next 	=(refr_tick && mushroom_stage_reg==6) ?(wall_y_t+3)// 6: begin
				: (refr_tick && mushroom_stage_reg==7) ? 479 				//7 : disappear
				: (refr_tick && mushroom_stage_reg==3) ? (mushroom_y_reg - 1)//3: up
				: (refr_tick && mushroom_stage_reg==4) ? (mushroom_y_reg + 4)//4: down
				: (refr_tick && mushroom_stage_reg==5) ? ( GROUND_Y_T - mushroom_hi_size) //5: back to base
				: (mushroom_y_reg);	
	assign mushroom_stage_next=((mario_x_l<=mushroom_x_r)&&(mario_x_l >= mushroom_x_l-mario_lo_size)&&(mario_y_t <= mushroom_y_b)&&(mario_y_t>=mushroom_y_t-mario_hi_size))? 7 // disappear
							:(mushroom_x_l <=6||mushroom_stage_reg==7) ? 				7 // disappear
							:(mushroom_x_r >= pipe1_x_l||mushroom_stage_reg==2)? 		2 // left
							:(mushroom_y_t == GROUND_Y_T-mushroom_hi_size)?		1 // right 
							:(mushroom_y_t > GROUND_Y_T-mushroom_hi_size)?		5 // back to base
							:(mushroom_x_l >= wall_x_r) ? 		4	// down
							:(mushroom_y_t <= wall_y_t -mushroom_hi_size) ?  	1	// right
							:((mario_x_l>=wall_x_l+25)&&(mario_x_l<=wall_x_l+50)&&(mario_y_t <=wall_y_b+6)&&(mario_y_t >= wall_y_b-6)&&(mushroom_stage_reg==6)) ? 3	//up
							: mushroom_stage_reg;

	//--------------------------DRAW MUSHROOM--------1-----------------------------------
	wire [4:0] rom_addr_mus;
	wire [4:0] rom_col_mus;
	reg [29:0] rom_data_mus;
	wire rom_bit_mus;
	wire rd_mus_on;	
	
	always @*
	case(rom_addr_mus)

		5'd0 :  rom_data_mus =  25'b0000000000000000000000000;
		5'd1 :  rom_data_mus =  25'b0000000000011110000000000;
		5'd2 :  rom_data_mus =  25'b0000000001111111000000000;
		5'd3 :  rom_data_mus =  25'b0000000011111100100000000;
		5'd4 :  rom_data_mus =  25'b0000001111110000011000000;
		5'd5 :  rom_data_mus =  25'b0000001111110000001000000;
		5'd6 :  rom_data_mus =  25'b0000011111110000000100000;
		5'd7 :  rom_data_mus =  25'b0000111111111000000010000;
		5'd8 :  rom_data_mus =  25'b0000111111111100000110000;
		5'd9 :  rom_data_mus =  25'b0011000000111111111111100;
		5'd10 :  rom_data_mus = 25'b0011000000011111111111100;
		5'd11 :  rom_data_mus = 25'b0111000000011111111001100;
		5'd12 :  rom_data_mus = 25'b0110000000001111111000110;
		5'd13 :  rom_data_mus = 25'b0110000000001111110000010;
		5'd14 :  rom_data_mus = 25'b0111000000011111111000010;
		5'd15 :  rom_data_mus = 25'b0111100000111111111100110;
		5'd16 :  rom_data_mus = 25'b0011111111111111111111100;
		5'd17 :  rom_data_mus = 25'b0000000011111111100000000;
		5'd18 :  rom_data_mus = 25'b0000000001111111000000000;
		5'd19 :  rom_data_mus = 25'b0000000011111111100000000;
		5'd20 :  rom_data_mus = 25'b0000000011111111100000000;
		5'd21 :  rom_data_mus = 25'b0000000011111111100000000;
		5'd22 :  rom_data_mus = 25'b0000000011111111100000000;
		5'd23 :  rom_data_mus = 25'b0000000001111111000000000;
		5'd24 :  rom_data_mus = 25'b0000000000000000000000000;
	endcase
	
	assign rom_addr_mus  = pix_y [4:0] - mushroom_y_t[4:0] ; //3bits
	assign rom_col_mus  = pix_x [4:0] - mushroom_x_l[4:0] ; //1 bit
	assign rom_bit_mus = rom_data_mus [rom_col_mus] ; 
	assign rd_mus_on  = sq_mushroom_on & rom_bit_mus;
				
	
	//--------------------------DRAW DRAGON--------1-----------------------------------
	wire [6:0] rom_addr_d;
	wire [6:0] rom_col_d;
	reg [75:0] rom_data_d;
	wire rom_bit_d;
	wire rd_d_on;	
	
	always @*
	case(rom_addr_d)

			7'd0 :  rom_data_d = 76'b0000000000000000000000000000000110111100000000000000000000000000000000000000;
			7'd1 :  rom_data_d = 76'b0000000000000000000000000000000010001000000000000000000000000000000000000000;
			7'd2 :  rom_data_d = 76'b0000000000000000000001100000001101101101110000000000000000000000000000000000;
			7'd3 :  rom_data_d = 76'b0000000000000000000111000000111111110100111100000000000000000000000000000000;
			7'd4 :  rom_data_d = 76'b0000000000000000011110000000111111011010001111000000000000000000000000000000;
			7'd5 :  rom_data_d = 76'b0000000000000011110110000000111111001111001001100000000000000000000000000000;
			7'd6:   rom_data_d = 76'b0000000000001111100100000000011100000101110000111000000000000000000000000000;
			7'd7 :  rom_data_d = 76'b0000000000000000001101100100000000000111000001010000000111000000000000000000;
			7'd8 :  rom_data_d = 76'b0000000000000000111001001100000001111111000000100001110011100000000000000000;
			7'd9 :  rom_data_d = 76'b0000000000000011100001111000000011011101100000110110011000110000000000000000;
			7'd10 : rom_data_d = 76'b0000000000000111001000011000001100001111110000011111001100011000000000000000;
			7'd11:  rom_data_d = 76'b0000000000011100011100011000011001111111110010001101100110001000000000000000;
			7'd12 : rom_data_d = 76'b0000000000111001110110010000010111001011111011001100101011001110000000000000;
			7'd13 : rom_data_d = 76'b0000000001100011000010010000101111011111011001000110111100100010000000000000;
			7'd14 : rom_data_d = 76'b0000000011000110000010100000101101111100101001100010011011011001000000000000;
			7'd15 : rom_data_d = 76'b0000000110001111101100100000011111111111111100110001010001111001110000000000;
			7'd16 : rom_data_d = 76'b0000001100011010111110100001110011100011101110110001001000111100011000000000;
			7'd17 : rom_data_d = 76'b0000001100110100010010000001111111100111011011111001101000011111001100000000;
			7'd18 : rom_data_d = 76'b0000011000101101100010010000100111000110001111111001101100001111000100000000;
			7'd19 : rom_data_d = 76'b0000011001011000100111110000111011000001100111110110000100000011100110000000;
			7'd20 : rom_data_d = 76'b0000000011110011000011000001101111100000011110111110000000000001110001000000;
			7'd21 : rom_data_d = 76'b0000010010100011000011000001100011111000001111111100000000000000111001000000;
			7'd22 : rom_data_d = 76'b0000110111100011000011011001111111011000000111101110000000000000011001100000;
			7'd23 : rom_data_d = 76'b0000101101000000000000111011100111000000001111111011100000000000010100110000;
			7'd24 : rom_data_d = 76'b0000100110000000000000101111111111101100001111110100000110000000001110110000;
			7'd25 : rom_data_d = 76'b0001101010000000000011010110111111101100010111110100001111000000001110010000;
			7'd26 : rom_data_d = 76'b0001011100000000000001011000111101011100110001110001111111110000000110010000;
			7'd27 : rom_data_d = 76'b0001011100000000000000111100000001011111000000000111111101111011000011011000;
			7'd28 : rom_data_d = 76'b0011011000000000000000001111000110000111100111111110110010111111000011011000;
			7'd29 : rom_data_d = 76'b0000111000000000000000010110001100100111111100001110110001001111100001101100;
			7'd30 : rom_data_d = 76'b0010011000000000000000010110011000110110011000000110010000101011010001101000;
			7'd31 : rom_data_d = 76'b0010110000000000000011101110010001010110011000001100011111011111011001110100;
			7'd32 : rom_data_d = 76'b0100100000000000000111111010100110110110001111111110111011111010001000100100;
			7'd33 : rom_data_d = 76'b0111110000011100001101110011111101101101100011000011110001001011000100110000;
			7'd34 : rom_data_d = 76'b0111100000011000011001110011110110001001110010000011111000110011000010111000;
			7'd35 : rom_data_d = 76'b0000100000110000010001100010001100111101011110001110011000010011000010011110;
			7'd36 : rom_data_d = 76'b0011100000100000110011000110110001111001101100011111111010001011000001001110;
			7'd37 : rom_data_d = 76'b0111000001000001100011000100111011110011000111001111111111110011000001101000;
			7'd38 : rom_data_d = 76'b1101000001100001000010011101111111000111000010110110010101111110000000101100;
			7'd39 : rom_data_d = 76'b1101100010111001000000110011001010001110000100110110011111111111000000101100;
			7'd40 : rom_data_d = 76'b1101100011111110001111111010001100111100011101110111111111111111111000010110;
			7'd41 : rom_data_d = 76'b1101100111001111111110000110001111110001111111010110000000001001111100011111;
			7'd42 : rom_data_d = 76'b0001101111110110111000001100010011100011100011110011100000000000000000001011;
			7'd43 : rom_data_d = 76'b0001111110100110001000001111110011000111000110110111101000000000000000001011;
			7'd44 : rom_data_d = 76'b0111101111100110001111100110111011111100011100111000111000000000000000000111;
			7'd45 : rom_data_d = 76'b0111100111011111111100011000101100011000111001110001111100000000000000000011;
			7'd46 : rom_data_d = 76'b0001001001111001111000000001101100111111100011000001101000000000000000000011;
			7'd47 : rom_data_d = 76'b0011101011000000011000000000101001110111000110000000110000000000000000000011;
			7'd48 : rom_data_d = 76'b0011101010000000110000000011111011100111111100110000111000000000000000000011;
			7'd49 : rom_data_d = 76'b0001101000000000100000000011011011000110111001110000001100000000000000000011;
			7'd50 : rom_data_d = 76'b0011010000000000000000000011011001000110111111100000001000000000000000000000;
			7'd51 : rom_data_d = 76'b0001110000000000000000000000010010000111011111000000000000000000000000000000;
			7'd52 : rom_data_d = 76'b0001100000000000000000000001111010000110010111100000100100000000000000000000;
			7'd53 : rom_data_d = 76'b0000110000000000000000000001001000001111111101100000110100000000000000000000;
			7'd54 : rom_data_d = 76'b0000111100000000000000000001101100011111111000000000111100000000000000000000;
			7'd55 : rom_data_d = 76'b0000011100000000000000000001111110001110010000100000110000000000000000000000;
			7'd56 : rom_data_d = 76'b0000011100000000000000000000100011111100100001100000100110000000000000000000;
			7'd57 : rom_data_d = 76'b0000001100000000000000000000110111111101100111010001100110000000000000000000;
			7'd58 : rom_data_d = 76'b0000001100000000000000000000010110101101101110001111000010000000000000000000;
			7'd59 : rom_data_d = 76'b0000000110000000000000000000001100111001110011001100011110000000000000000000;
			7'd60 : rom_data_d = 76'b0000000000000000000000000000000111011111000001111111111110000000000000000000;
			7'd61 : rom_data_d = 76'b0000000000000000000000000000000011011010010000110111110010000000000000000000;
			7'd62 : rom_data_d = 76'b0000000000000000000000000000000000011010001011100110010000000000000000000000;
			7'd63 : rom_data_d = 76'b0000000000000000000000000000000001011111111110000000000000000000000000000000;
			7'd64 : rom_data_d = 76'b0000000000000000000000000000000011000001110000000000011010000000000000000000;
			7'd65 : rom_data_d = 76'b0000000000000000000000000000000011010000000000000000001010000000000000000000;
			7'd66 : rom_data_d = 76'b0000000000000000000000000000000010111100000000000111011111000000000000000000;
			7'd67 : rom_data_d = 76'b0000000000000000000000000000000010101100000000000111010111000000000000000000;
			7'd68 : rom_data_d = 76'b0000000000000000000000000000000000001100000000000001110010000000000000000000;
			7'd69 : rom_data_d = 76'b0000000000000000000000000000000000000000000000000010110011000000000000000000;
			7'd70 : rom_data_d = 76'b0000000000000000000000000000000000000000000000000010010000000000000000000000;
		endcase
	
	
	//-----------------------------DRAW DRAGON -----------------------------	
	
	assign rom_addr_d  = pix_y [6:0] - monster_y_t[6:0] ; //3bits
	assign rom_col_d  = pix_x [6:0] - monster_x_l[6:0] ; //1 bit
	assign rom_bit_d  = rom_data_d [rom_col_d] ; 
	assign rd_d_on  = monster_on & rom_bit_d;	
	
	
	
	//----------------------Turn on 
	// use to built sence for game
	reg pipe1_turn_next, pipe1_turn_reg;
	reg pri_turn_next, pri_turn_reg;
	reg wall_turn_next, wall_turn_reg;

	reg hole1_turn_next, hole1_turn_reg;
	reg turn_again;
	
	always@*
	if(refr_tick)
		begin

			pipe1_turn_next = 1;

			wall_turn_next = wall_turn_reg;
			hole1_turn_next = hole1_turn_reg;

			wall_lo_size_next = wall_lo_size_reg;
			wall_y_next <= wall_y_reg;
			
				begin
					//--------------------------------- scene 1
					if (built_reg == 0 ) begin wall_turn_next = 1; wall_y_next <=300; wall_lo_size_next <= mario_lo_size * 6 ; end//  wall appear at beginning			
					else if(wall_x_l <= 1 )	begin	wall_turn_next = 0; end

					//--------------------------------- scene 2					
					//165 is time that object appear again
					if (built_reg == 165 ) begin wall_turn_next = 1; wall_y_next <= 300;  wall_lo_size_next <= 200;end					
					else if(wall_x_l <= 1 )	begin	wall_turn_next = 0;  end
					
					if (built_reg == 135 ) begin hole1_turn_next = 1; end //hole appear
					else if(hole1_x_l <= 1 )	begin	hole1_turn_next = 0;  end					
				end				
		end	
	
		//------------------------------- MARIO DEAD
	reg dead_next, dead_reg;
	
	always@*
	begin
		dead_next = dead_reg;
		//update mario dead when he drop the the hole
		if (mario_y_t >= MAX_Y)  dead_next = 1; 
		
		//update mario dead when he touch Dragon
		else if((mario_x_l<=mushroom_x_r)&&(mario_x_l >= mushroom_x_l-mario_lo_size)&&(mario_y_t <= mushroom_y_b)&&(mario_y_t>=mushroom_y_t-mario_hi_size))
			begin big_next=1;shift=1;end
		else if ( mst_turn_reg && (monster_x_l - mario_lo_size + 1 < mario_x_l) && (mario_x_l < monster_x_r - 1) 
               &&  (monster_y_t - 1 < mario_y_t) && (mario_y_t < monster_y_b - 1))
            if(big)
				begin big_next=0;shift=1;end
			else
				dead_next = 1;
		//update mario dead when he touch Goompa(small monster)
		else if (goo_turn_reg && (goo_x_l - mario_lo_size + 1 < mario_x_l) && (mario_x_l < goo_x_r - 1) 
               &&  (goo_y_t +4 < mario_y_b) && (mario_y_t < goo_y_b - 1))
		    if(big)
				begin big_next=0;shift=1;end
			else
				dead_next = 1;
		else if(~KEY[3] & ~KEY[2])  dead_next = 0; //press both key to reset game 
		else
			begin  big_next=big;shift=0;end
	end	
	
	
	//update the mario dead
	always@(posedge CLOCK_50)
		begin
			dead_reg <= dead_next;
		end
	//------------------------------- DRAGON DEAD
	always@*
		begin
			//update for Dragon
			goo_turn_next =goo_turn_reg;
			mst_turn_next = mst_turn_reg;
			pri_turn_next=pri_turn_reg;
			if (built_reg == 165 ) mst_turn_next = 1;// Dragon appear
			else if((monster_y_t + 10 > mario_y_b) && (monster_y_t - 10 < mario_y_b) 
					&& (monster_x_l < mario_x_l) && (monster_x_r > mario_x_r)) begin mst_turn_next = 0;pri_turn_next =1;end // dragon dead when mario is on his head
					
			//update for goompa dead
			if (built_reg == 165 ) goo_turn_next = 1;//Goopa appear
			else 
					if((goo_y_t + 4 > mario_y_b) && (goo_y_t - 4 < mario_y_b)
					&& ((goo_x_l <= mario_x_l) && (goo_x_r > mario_x_r )
					|| (goo_x_l >= mario_x_l) && (goo_x_l <= mario_x_r + 3)
					|| (goo_x_r > mario_x_l + 3) && (goo_x_r <= mario_x_r)))
					 goo_turn_next = 0;		//goompa dead when mario in on his head
					
		end	
	
	
    //--------------------------------------------GOOMPA----------------------------------------------
	localparam GOO_X = 30;
	localparam GOO_Y = 29;
	reg goo_turn_reg;
    reg goo_turn_next;
	wire [9:0] goo_x_l, goo_x_r, goo_y_t, goo_y_b;
	reg [9:0] goo_x_reg, goo_y_reg;
	wire [9:0] goo_x_next, goo_y_next;
	reg  [9:0] gooX_delta_reg ,gooX_delta_next ; 
	reg  [9:0] gooY_delta_reg, gooY_delta_next;
	localparam  GOO_V_P = 2;
	localparam  GOO_V_N = -2; 
	wire goo_on;
	wire [8:0] goo_rgb;
	
	
	//--------------------------DRAW GOOMPA--------1-----------------------------------
	wire [4:0] rom_addr_goo;
	wire [4:0] rom_col_goo;
	reg [29:0] rom_data_goo;
	wire rom_bit_goo;
	wire rd_goo_on;
	
	
	always @*
	case(rom_addr_goo)

		5'd0 :  rom_data_goo =  30'b000000000000000000000000000000;
		5'd1 :  rom_data_goo =  30'b000000000000111111100000000000;
		5'd2 :  rom_data_goo =  30'b000000000000111111100000000000;
		5'd3 :  rom_data_goo =  30'b000000000011111111111000000000;
		5'd4 :  rom_data_goo =  30'b000000001111111111111110000000;
		5'd5 :  rom_data_goo =  30'b000000001111111111111110000000;
		5'd6 :  rom_data_goo =  30'b000000111111111111111111100000;
		5'd7 :  rom_data_goo =  30'b000000111111111111111111100000;
		5'd8 :  rom_data_goo =  30'b000011111111111111111111111000;
		5'd9 :  rom_data_goo =  30'b000011111111111111111111111000;
		5'd10 :  rom_data_goo = 30'b001111111011111111111001111100;
		5'd11 :  rom_data_goo = 30'b001111110011111111111001111110;
		5'd12 :  rom_data_goo = 30'b001111110011111111111001111100;
		5'd13 :  rom_data_goo = 30'b111111110011111111111001111111;
		5'd14 :  rom_data_goo = 30'b111111110011001110011001111111;
		5'd15 :  rom_data_goo = 30'b111111110011001111011001111111;
		5'd16 :  rom_data_goo = 30'b111111110000001111000001111111;
		5'd17 :  rom_data_goo = 30'b111111111111111111111111111111;
		5'd18 :  rom_data_goo = 30'b111111111111111111111111111111;
		5'd19 :  rom_data_goo = 30'b001111111100000000000111111110;
		5'd20 :  rom_data_goo = 30'b001111110000000000000001111100;
		5'd21 :  rom_data_goo = 30'b000000000000000000000001000000;
		5'd22 :  rom_data_goo = 30'b000011110000000000000001000000;
		5'd23 :  rom_data_goo = 30'b000011111000000000000000000000;
		5'd24 :  rom_data_goo = 30'b001111111111000000000111100000;
		5'd25 :  rom_data_goo = 30'b001111111111100000001111100000;
		5'd26 :  rom_data_goo = 30'b011111111111110000011111110000;
		5'd27 :  rom_data_goo = 30'b000111111111111100111111111100;
		5'd28 :  rom_data_goo = 30'b000001111111111111111111111100;
	endcase
					
		assign rom_addr_goo  = pix_y [4:0] - goo_y_t[4:0] ; //3bits
		assign rom_col_goo  = pix_x [4:0] - goo_x_l[4:0] ; //1 bit
		assign rom_bit_goo  = rom_data_goo [rom_col_goo] ; 
		assign rd_goo_on  = goo_on & rom_bit_goo;
	

	// ----------Registers---------------
	always@(posedge CLOCK_50,posedge reset, posedge dead_reg)
		if(reset  | dead_reg)	
			begin
				vr = 10'h002;			
				max_jump = 150;
				Drop_reg <= 0;
				state_reg <= 2;
				at_mid_reg <= 0;			
				//vr <= 10'h002;
				mario_base_reg <= BASE;
				
				mario_x_reg <= 100;      //initial position x mario
				mario_y_reg <= 385;
				big <=0;
				mario_del_run_reg <= 10'h002;
				mario_del_jump_reg <= 10'h002;
				mario_highest_reg <= mario_base_reg - max_jump;			
				//wall_x_del_reg <= 0;  
				wall_x_reg <= 369;        //wall initial at  high is constant
				pipe1_x_reg <= 639;
				hole1_x_reg <= 639;
				c_x_reg <= 100;
				c1_x_reg <= 400;
				//Built Counter
				built_reg <= 0;
				wall_turn_reg <= 1;
				pipe1_turn_reg <= 0;
				hole1_turn_reg <= 0;
				
								
				//monster
				mst_turn_reg <= 0;
				monster_x_reg <= MAX_X;
				monster_y_reg <= 0;				
				mstX_delta_reg <= 5;
				mstY_delta_reg <= 5;
				
				//goompa
				goo_turn_reg <= 1;
				goo_x_reg <= 639;
				goo_y_reg <= GROUND_Y_T;		
				gooX_delta_reg <= 5;
				gooY_delta_reg <= 5;
				//mushroom
				mushroom_stage_reg <= 6; // begin
				mushroom_x_reg <= wall_x_l+25;
				mushroom_y_reg <= wall_y_t;
				pri_turn_reg <=0;
				pri_x_reg <= 639;
			end
		else
			begin
				pri_turn_reg <= pri_turn_next;
				pri_x_reg <= pri_x_next;
				vr = vr_next;
				max_jump = max_jump_next;
				Drop_reg <= Drop_next;
				state_reg <= state_next;
				at_mid_reg <= at_mid_next;
				//Built counter
				built_reg <= built_next;				
				//Turn on
				wall_turn_reg <= wall_turn_next;
				pipe1_turn_reg <= pipe1_turn_next;
				hole1_turn_reg <= hole1_turn_next;				
				
				//--------------MONSTER
				monster_x_reg <= monster_x_next;
				monster_y_reg <= monster_y_next;
				mstX_delta_reg <= mstX_delta_next; 
				mstY_delta_reg <= mstY_delta_next;
				mst_turn_reg <= mst_turn_next;
				
				//--------------GOOPA CLOCK
				goo_x_reg <= goo_x_next;
				goo_y_reg <= goo_y_next;
				gooX_delta_reg <=gooX_delta_next; 
				gooY_delta_reg <=gooY_delta_next;
				goo_turn_reg <=goo_turn_next;
				
				//--------------MARIO
				mario_del_run_reg = mario_del_run_next;
				mario_del_jump_reg = mario_del_jump_next;				
				mario_base_reg = mario_base_next;
				mario_highest_reg <= mario_highest_next;				
				mario_x_reg <= mario_x_next;
				mario_y_reg <= mario_y_next;
				big = big_next;
				
				//positon of objects
				wall_lo_size_reg <= wall_lo_size_next; // change at built
				wall_x_reg <= wall_x_next;
				wall_y_reg <= wall_y_next; // change at built
				
				//pipe1  hole   cloud
				pipe1_x_reg <= pipe1_x_next;				
				hole1_x_reg <= hole1_x_next;
				c_x_reg <= c_x_next;
				c1_x_reg <= c1_x_next;
				//mushroom
				mushroom_stage_reg=mushroom_stage_next;
				mushroom_x_reg=mushroom_x_next;
				mushroom_y_reg=mushroom_y_next;	
			end

		assign refr_tick = (pix_x == 0) && (pix_y == 481);
		assign at_mid_next = (mario_x_reg >= (MAX_X) /2 - 30 ) ? 1 : 0;
		
		//Built counter		
		assign built_next = (refr_tick & at_mid_reg & slo_clk & mario_del_run_next != 0) ? built_reg + 1 : built_reg;	
		reg [5:0]vir_clk = 0;
		reg slo_clk;
		always@(posedge refr_tick)
			begin
				vir_clk = vir_clk + 1;
				slo_clk = vir_clk[3];
			end
			
			
		//update the highest level that mario can jump to
		always@*
			if(big)
				max_jump_next =  150 + 64 ; // mario can jump higher when he big
			else  
				max_jump_next =  150;
				
			//-----------------------------GROUND-----------------------------
		assign ground_on = (GROUND_Y_T <= pix_y) && (pix_y <= GROUND_Y_B); 
			
			//-------------------------------MONSTER--------------------------------
		localparam monster_hi_max = 430;
		localparam monster_lo_max = 600;
		assign monster_x_l = monster_x_reg;
		assign monster_x_r = monster_x_l + MONSTER_X - 1;		 
		assign monster_y_b = monster_y_reg;      		                                   
		assign monster_y_t = monster_y_b - MONSTER_Y - 1;
		assign monster_on = (monster_x_l <= pix_x) && (pix_x <= monster_x_r) && (monster_y_t <= pix_y) && (pix_y <= monster_y_b);
		assign monster_rgb = 9'b0;//black color

		assign monster_x_next  =  (mst_turn_reg) & (refr_tick)  ?  monster_x_reg + mstX_delta_reg  : monster_x_reg;  
		assign monster_y_next  =  (mst_turn_reg & refr_tick)  ?  monster_y_reg + mstY_delta_reg  : monster_y_reg;
		//update moving for Monster
		always @*
			if(mst_turn_reg)
			begin		
			 mstY_delta_next = mstY_delta_reg;
			 mstX_delta_next = mstX_delta_reg;
			 if(monster_y_t < 100)
			     mstY_delta_next = MONSTER_V_P;
			 else if(monster_y_b > monster_hi_max)
			     mstY_delta_next = MONSTER_V_N;
			 else if (monster_x_l < 1)
			     mstX_delta_next = MONSTER_V_P;
			 else if (monster_x_r > monster_lo_max)
			     mstX_delta_next = MONSTER_V_N;
		end

		//-------------------------GOOMPA-------------------------------------
		localparam goo_hi_max = 430;
		localparam goo_lo_max = 600;
		assign goo_x_l = goo_x_reg;
		assign goo_x_r = goo_x_l + GOO_X - 1;		 
		assign goo_y_b = goo_y_reg;      		                                   
		assign goo_y_t = goo_y_b - GOO_Y - 1;
		assign goo_on = (goo_x_l <= pix_x) && (pix_x <= goo_x_r) && (goo_y_t <= pix_y) && (pix_y <= goo_y_b);
		assign goo_rgb = 9'b0;

		assign goo_x_next  =  (goo_turn_reg) & (refr_tick)  ?  goo_x_reg + gooX_delta_reg  : goo_x_reg;  
		assign goo_y_next  =  (goo_turn_reg & refr_tick)  ?  goo_y_reg  : goo_y_reg;

		//update position (moving) of goompa (small monster)
		always @*
			if(goo_turn_reg)
			begin			
				gooY_delta_next =gooY_delta_reg;
				gooX_delta_next =gooX_delta_reg;
				 if (goo_x_l < 3)
					gooX_delta_next = GOO_V_P;
				 else if (goo_x_r > goo_lo_max)
					gooX_delta_next = GOO_V_N;
			end
		
		
	//-----------------------------CLOUD-----------------------------
			
		assign c_x_l = c_x_reg;
		assign c_y_t = 100;
		assign c_x_r  = c_x_l  + C_LO_SIZE - 1;
		assign c_y_b  = c_y_t  + C_HI_SIZE - 1; 
		assign sq_c_on = (c_x_l <= pix_x) && (pix_x <= c_x_r) && (c_y_t <= pix_y)  && (pix_y <= c_y_b);
		//draw cloud
		assign rom_addr_c  = pix_y [3:0] - c_y_t[3:0] ; //3bits
		assign rom_col_c  = pix_x [5:0] - c_x_l[5:0] ; //1 bit
		assign rom_bit_c  = rom_data_c [rom_col_c] ; 
		assign rd_c_on  = sq_c_on & rom_bit_c;
		
		//update the positon of cloud
		always@*			
			begin
				c_x_next = c_x_reg;
				if(refr_tick & ~KEY[0] & at_mid_reg )
					c_x_next = c_x_reg - mario_del_run_next;
			end
		
		
		
		//----------------- WALL--------------------------------------		
		assign rom_addr_w  = pix_y [4:0] - wall_y_t[4:0] ; //3bits
		assign rom_col_w  = pix_x [7:0] - wall_x_l[7:0] ; //1 bit
		assign rom_bit_wall  = rom_data_w [rom_col_w] ; 
		assign rd_wall_on  = wall_on & rom_bit_wall;   
  
		assign wall_y_t = wall_y_reg;
		assign wall_x_l = wall_x_reg;
		assign wall_y_b = wall_y_t + wall_hi_size - 1;
		assign wall_x_r = wall_x_l + wall_lo_size_reg - 1;
		assign wall_on = ( wall_x_l <= pix_x ) && (pix_x <= wall_x_r) && (wall_y_t <= pix_y) && (pix_y <= wall_y_b)  ;
		
		//update the postion of wall
		always@*			
			begin				
				wall_x_next = wall_x_reg;
				if (built_reg == 165 ) wall_x_next = 639;//wall appear again at built_reg == 165
				else if(wall_turn_reg & refr_tick & ~KEY[0] & at_mid_reg )
					wall_x_next = wall_x_reg - mario_del_run_next;
			end
		
		
		
		//----------------PIPE1-----------------------------------------			
		assign pipe1_y_b = pipe1_y_t + pipe1_hi_size - 1;
		assign pipe1_x_l = pipe1_x_reg;
		assign pipe1_x_r = pipe1_x_l + pipe1_lo_size - 1;	
		assign rd_pipe1_on = ( pipe1_x_l <= pix_x ) && (pix_x <= pipe1_x_r) && (pipe1_y_t <= pix_y) && (pix_y <= pipe1_y_b);
			
		//update the position of base			
		always@*			
			begin
				pipe1_x_next = pipe1_x_reg;
				if( pipe1_turn_reg & refr_tick & ~KEY[0] & at_mid_reg)					
					pipe1_x_next = pipe1_x_reg - mario_del_run_next;					
			end
			
		
		//----------------HOLE1-----------------------------------------
		assign hole1_y_t = BASE;
		assign hole1_y_b = hole1_y_t + hole1_hi_size - 1;
		assign hole1_x_l = hole1_x_reg;
		assign hole1_x_r = hole1_x_l + hole1_lo_size - 1;
		
		assign hole1_on = ( hole1_x_l <= pix_x ) && (pix_x <= hole1_x_r) && (hole1_y_t <= pix_y) && (pix_y <= hole1_y_b);			
		assign hole1_rgb = backgroud_rgb;				
		
		//update moving of hole1
		always@*			
			begin
				hole1_x_next = hole1_x_reg;
				if (built_reg == 135) hole1_x_next = 639; //this code is to call the hole appear again at time built_reg == 135
				else if( hole1_turn_reg & refr_tick & ~KEY[0] & at_mid_reg)					
					hole1_x_next = hole1_x_reg - mario_del_run_next;
		end
		
		//-------------------------BEGIN MARIO--------------------------------------------------------------------------------------------------


		assign mario_x_l = mario_x_reg;
		assign mario_y_t = mario_y_reg;	
		assign mario_x_r = mario_x_l + mario_lo_size;
		assign mario_y_b = mario_y_t + mario_hi_size;

		reg red1,red2,red3,red4,red5,red6,red7,red8,red9,red10,red11;
		reg blue1,blue2,blue3,blue4,blue5,blue6,blue7,blue8,blue9,blue10;
		reg yellow1,yellow2,yellow3,yellow4,yellow5,yellow6,yellow7,yellow8,yellow9,yellow10,yellow11,yellow12,yellow13;
		reg black1,black2,black3,black4,black5,black6,black7,black8,black9,black10,black11,black12;
		wire mario_red,mario_blue,mario_yellow,mario_black;
		assign mario_red=red1||red2||red3||red4||red5||red6||red7||red8||red9||red10||red11;
		assign mario_blue=blue1||blue2||blue3||blue4||blue5||blue6||blue7||blue8||blue9||blue10;
		assign mario_yellow=yellow1||yellow2||yellow3||yellow4||yellow5||yellow6||yellow7||yellow8||yellow9||yellow10||yellow11||yellow12||yellow13;
		assign mario_black=black1||black2||black3||black4||black5||black6||black7||black8||black9||black10||black11||black12;
		always @*
		begin
		
		if(big)
		begin//draw the big mario
			mario_hi_size=64;
			mario_lo_size=36;
			
			red1=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 36) && (mario_y_t +4 <= pix_y) && (pix_y <= mario_y_t +8);
			red2=(mario_x_l +9 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t <= pix_y) && (pix_y <= mario_y_t +4);
			red3=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 12) && (mario_y_t +28 <= pix_y) && (pix_y <= mario_y_t +32);
			red4=(mario_x_l +15 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +28<= pix_y) && (pix_y <= mario_y_t +32);	
			red5=(mario_x_l +3 <= pix_x) && ( pix_x <= mario_x_l + 12) && (mario_y_t +32<= pix_y) && (pix_y <= mario_y_t +36);
			red6=(mario_x_l +15 <= pix_x) && ( pix_x <= mario_x_l + 21) && (mario_y_t +32<= pix_y) && (pix_y <= mario_y_t +36);
			red7=(mario_x_l +24 <= pix_x) && ( pix_x <= mario_x_l + 33) && (mario_y_t +32<= pix_y) && (pix_y <= mario_y_t +36);
			red8=(mario_x_l  <= pix_x) && ( pix_x <= mario_x_l + 12) && (mario_y_t +36<= pix_y) && (pix_y <= mario_y_t +40);
			red9=(mario_x_l +24 <= pix_x) && ( pix_x <= mario_x_l + 36) && (mario_y_t +36<= pix_y) && (pix_y <= mario_y_t +40);
			red10=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 9) && (mario_y_t +40<= pix_y) && (pix_y <= mario_y_t +44);
			red11=(mario_x_l +27 <= pix_x) && ( pix_x <= mario_x_l + 30) && (mario_y_t +40<= pix_y) && (pix_y <= mario_y_t +44);


			blue1=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 15) && (mario_y_t +52 <= pix_y) && (pix_y <= mario_y_t +56);
			blue2=(mario_x_l +21 <= pix_x) && ( pix_x <= mario_x_l + 30) && (mario_y_t +52 <= pix_y) && (pix_y <= mario_y_t +56);
			blue3=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 30) && (mario_y_t +48 <= pix_y) && (pix_y <= mario_y_t +52);
			blue4=(mario_x_l +9 <= pix_x) && ( pix_x <= mario_x_l + 27) && (mario_y_t +44 <= pix_y) && (pix_y <= mario_y_t +48);
			blue5=(mario_x_l +9 <= pix_x) && ( pix_x <= mario_x_l + 12) && (mario_y_t +40 <= pix_y) && (pix_y <= mario_y_t +44);
			blue6=(mario_x_l +15 <= pix_x) && ( pix_x <= mario_x_l + 21) && (mario_y_t +40 <= pix_y) && (pix_y <= mario_y_t +44);
			blue7=(mario_x_l +24 <= pix_x) && ( pix_x <= mario_x_l + 27) && (mario_y_t +40 <= pix_y) && (pix_y <= mario_y_t +44);
			blue8=(mario_x_l +21 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +36 <= pix_y) && (pix_y <= mario_y_t +40);
			blue9=(mario_x_l +12 <= pix_x) && ( pix_x <= mario_x_l + 15) && (mario_y_t +28 <= pix_y) && (pix_y <= mario_y_t +36);
			blue10=(mario_x_l +21 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +32 <= pix_y) && (pix_y <= mario_y_t +36);

			yellow1=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 9) && (mario_y_t +12 <= pix_y) && (pix_y <= mario_y_t +20);
			yellow2=(mario_x_l +12 <= pix_x) && ( pix_x <= mario_x_l + 15) && (mario_y_t +12 <= pix_y) && (pix_y <= mario_y_t +16);
			yellow3=(mario_x_l +9 <= pix_x) && ( pix_x <= mario_x_l + 21) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t +28);
			yellow4=(mario_x_l +21 <= pix_x) && ( pix_x <= mario_x_l + 30) && (mario_y_t +24 <= pix_y) && (pix_y <= mario_y_t +28);
			yellow5=(mario_x_l +15 <= pix_x) && ( pix_x <= mario_x_l + 21) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t +20);
			yellow6=(mario_x_l +21 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +16 <= pix_y) && (pix_y <= mario_y_t +20);
			yellow7=(mario_x_l +16 <= pix_x) && ( pix_x <= mario_x_l + 27) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t +16);
			yellow8=(mario_x_l +27 <= pix_x) && ( pix_x <= mario_x_l + 33) && (mario_y_t +12 <= pix_y) && (pix_y <= mario_y_t +20);
			yellow9=(mario_x_l +33 <= pix_x) && ( pix_x <= mario_x_l + 36) && (mario_y_t +16 <= pix_y) && (pix_y <= mario_y_t +20);
			yellow10=(mario_x_l  <= pix_x) && ( pix_x <= mario_x_l + 6) && (mario_y_t +40 <= pix_y) && (pix_y <= mario_y_t +52);
			yellow11=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 9) && (mario_y_t +44 <= pix_y) && (pix_y <= mario_y_t +48);
			yellow12=(mario_x_l +27 <= pix_x) && ( pix_x <= mario_x_l + 30) && (mario_y_t +44 <= pix_y) && (pix_y <= mario_y_t +48);
			yellow13=(mario_x_l +30  <= pix_x) && ( pix_x <= mario_x_l + 36) && (mario_y_t +40 <= pix_y) && (pix_y <= mario_y_t +52);

			black1=(mario_x_l +3 <= pix_x) && ( pix_x <= mario_x_l + 6) && (mario_y_t +12 <= pix_y) && (pix_y <= mario_y_t +24);
			black2=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 9) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t +24);
			black3=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 15) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t +12);
			black4=(mario_x_l +9 <= pix_x) && ( pix_x <= mario_x_l + 12) && (mario_y_t +12 <= pix_y) && (pix_y <= mario_y_t + 20);
			black5=(mario_x_l +12 <= pix_x) && ( pix_x <= mario_x_l + 15) && (mario_y_t +16 <= pix_y) && (pix_y <= mario_y_t + 20);
			black6=(mario_x_l +21 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t + 16);
			black7=(mario_x_l +24 <= pix_x) && ( pix_x <= mario_x_l + 27) && (mario_y_t +16 <= pix_y) && (pix_y <= mario_y_t + 20);
			black8=(mario_x_l +21 <= pix_x) && ( pix_x <= mario_x_l + 33) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t + 24);
			black9=(mario_x_l +0 <= pix_x) && ( pix_x <= mario_x_l + 3) && (mario_y_t +60 <= pix_y) && (pix_y <= mario_y_t + 64);
			black10=(mario_x_l +3 <= pix_x) && ( pix_x <= mario_x_l + 12) && (mario_y_t +56 <= pix_y) && (pix_y <= mario_y_t + 64);
			black11=(mario_x_l +24 <= pix_x) && ( pix_x <= mario_x_l + 33) && (mario_y_t +56 <= pix_y) && (pix_y <= mario_y_t + 64);
			black12=(mario_x_l +33 <= pix_x) && ( pix_x <= mario_x_l + 36) && (mario_y_t +60 <= pix_y) && (pix_y <= mario_y_t + 64);
		end
	
		else //Draw the small mario
		begin
			mario_hi_size=32;
			mario_lo_size=24;
			red1=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +2 <= pix_y) && (pix_y <= mario_y_t +4);
			red2=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 16) && (mario_y_t <= pix_y) && (pix_y <= mario_y_t +2);
			 red3=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 8) && (mario_y_t +14 <= pix_y) && (pix_y <= mario_y_t +16);
			 red4=(mario_x_l +10 <= pix_x) && ( pix_x <= mario_x_l + 16) && (mario_y_t +14<= pix_y) && (pix_y <= mario_y_t +16);	
			 red5=(mario_x_l +2 <= pix_x) && ( pix_x <= mario_x_l + 8) && (mario_y_t +16<= pix_y) && (pix_y <= mario_y_t +18);
			 red6=(mario_x_l +10 <= pix_x) && ( pix_x <= mario_x_l + 14) && (mario_y_t +16<= pix_y) && (pix_y <= mario_y_t +18);
			 red7=(mario_x_l +16 <= pix_x) && ( pix_x <= mario_x_l + 22) && (mario_y_t +16<= pix_y) && (pix_y <= mario_y_t +18);
			 red8=(mario_x_l  <= pix_x) && ( pix_x <= mario_x_l + 8) && (mario_y_t +18<= pix_y) && (pix_y <= mario_y_t +20);
			 red9=(mario_x_l +16 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +18<= pix_y) && (pix_y <= mario_y_t +20);
			 red10=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 6) && (mario_y_t +20<= pix_y) && (pix_y <= mario_y_t +22);
			 red11=(mario_x_l +18 <= pix_x) && ( pix_x <= mario_x_l + 20) && (mario_y_t +20<= pix_y) && (pix_y <= mario_y_t +22);


			 blue1=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 10) && (mario_y_t +26 <= pix_y) && (pix_y <= mario_y_t +28);
			 blue2=(mario_x_l +14 <= pix_x) && ( pix_x <= mario_x_l + 20) && (mario_y_t +26 <= pix_y) && (pix_y <= mario_y_t +28);
			 blue3=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 20) && (mario_y_t +24 <= pix_y) && (pix_y <= mario_y_t +26);
			 blue4=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 18) && (mario_y_t +22 <= pix_y) && (pix_y <= mario_y_t +24);
			 blue5=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 8) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t +22);
			 blue6=(mario_x_l +10 <= pix_x) && ( pix_x <= mario_x_l + 14) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t +22);
			 blue7=(mario_x_l +16 <= pix_x) && ( pix_x <= mario_x_l + 18) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t +22);
			 blue8=(mario_x_l +8 <= pix_x) && ( pix_x <= mario_x_l + 16) && (mario_y_t +18 <= pix_y) && (pix_y <= mario_y_t +20);
			 blue9=(mario_x_l +8 <= pix_x) && ( pix_x <= mario_x_l + 10) && (mario_y_t +14 <= pix_y) && (pix_y <= mario_y_t +18);
			 blue10=(mario_x_l +14 <= pix_x) && ( pix_x <= mario_x_l + 16) && (mario_y_t +16 <= pix_y) && (pix_y <= mario_y_t +18);

			 yellow1=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 6) && (mario_y_t +6 <= pix_y) && (pix_y <= mario_y_t +10);
			 yellow2=(mario_x_l +8 <= pix_x) && ( pix_x <= mario_x_l + 10) && (mario_y_t +6 <= pix_y) && (pix_y <= mario_y_t +8);
			 yellow3=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 14) && (mario_y_t +10 <= pix_y) && (pix_y <= mario_y_t +14);
			 yellow4=(mario_x_l +14 <= pix_x) && ( pix_x <= mario_x_l + 20) && (mario_y_t +12 <= pix_y) && (pix_y <= mario_y_t +14);
			 yellow5=(mario_x_l +10 <= pix_x) && ( pix_x <= mario_x_l + 14) && (mario_y_t +4 <= pix_y) && (pix_y <= mario_y_t +10);
			 yellow6=(mario_x_l +14 <= pix_x) && ( pix_x <= mario_x_l + 16) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t +10);
			 yellow7=(mario_x_l +16 <= pix_x) && ( pix_x <= mario_x_l + 18) && (mario_y_t +4 <= pix_y) && (pix_y <= mario_y_t +8);
			 yellow8=(mario_x_l +18 <= pix_x) && ( pix_x <= mario_x_l + 22) && (mario_y_t +6 <= pix_y) && (pix_y <= mario_y_t +10);
			 yellow9=(mario_x_l +22 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t +10);
			 yellow10=(mario_x_l  <= pix_x) && ( pix_x <= mario_x_l + 4) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t +26);
			 yellow11=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 6) && (mario_y_t +22 <= pix_y) && (pix_y <= mario_y_t +24);
			 yellow12=(mario_x_l +18 <= pix_x) && ( pix_x <= mario_x_l + 20) && (mario_y_t +22 <= pix_y) && (pix_y <= mario_y_t +24);
			 yellow13=(mario_x_l +20  <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +20 <= pix_y) && (pix_y <= mario_y_t +26);

			 black1=(mario_x_l +2 <= pix_x) && ( pix_x <= mario_x_l + 4) && (mario_y_t +6 <= pix_y) && (pix_y <= mario_y_t +12);
			 black2=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 6) && (mario_y_t +10 <= pix_y) && (pix_y <= mario_y_t +12);
			 black3=(mario_x_l +4 <= pix_x) && ( pix_x <= mario_x_l + 10) && (mario_y_t +4 <= pix_y) && (pix_y <= mario_y_t +6);
			black4=(mario_x_l +6 <= pix_x) && ( pix_x <= mario_x_l + 8) && (mario_y_t +6 <= pix_y) && (pix_y <= mario_y_t + 10);
			 black5=(mario_x_l +8 <= pix_x) && ( pix_x <= mario_x_l + 10) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t + 10);
			 black6=(mario_x_l +14 <= pix_x) && ( pix_x <= mario_x_l + 16) && (mario_y_t +4 <= pix_y) && (pix_y <= mario_y_t + 8);
			 black7=(mario_x_l +16 <= pix_x) && ( pix_x <= mario_x_l + 18) && (mario_y_t +8 <= pix_y) && (pix_y <= mario_y_t + 10);
			 black8=(mario_x_l +14 <= pix_x) && ( pix_x <= mario_x_l + 22) && (mario_y_t +10 <= pix_y) && (pix_y <= mario_y_t + 12);
			 black9=(mario_x_l  <= pix_x) && ( pix_x <= mario_x_l + 2) && (mario_y_t +30 <= pix_y) && (pix_y <= mario_y_t + 32);
			 black10=(mario_x_l +2 <= pix_x) && ( pix_x <= mario_x_l + 8) && (mario_y_t +28 <= pix_y) && (pix_y <= mario_y_t + 32);
			 black11=(mario_x_l +16 <= pix_x) && ( pix_x <= mario_x_l + 22) && (mario_y_t +28 <= pix_y) && (pix_y <= mario_y_t + 32);
			 black12=(mario_x_l +22 <= pix_x) && ( pix_x <= mario_x_l + 24) && (mario_y_t +30 <= pix_y) && (pix_y <= mario_y_t + 32);
		end
	end
		//update horizontal mario moving
		assign mario_x_next = (refr_tick && ~KEY[1]) ? (mario_x_reg - mario_del_run_next) //key[1]  is moving forward
							: (refr_tick && ~KEY[0] && ~at_mid_reg) ? (mario_x_reg + mario_del_run_next) //key[0] is moving backward
							: (mario_x_reg);
		//update vertical mario moving
		assign mario_y_next = (refr_tick && shift)? (mario_y_reg - 32) //shift the mario up with 32 pixel to prevent him stuck on ground when he eat mushroom
							:(refr_tick && state_reg == 0) ? (mario_y_reg  - mario_del_jump_reg) //up
							: (refr_tick && state_reg == 1) ? (mario_y_reg  + mario_del_jump_reg) //down
							: (refr_tick && state_reg == 2) ? (mario_y_reg) //no move
							:  mario_y_reg ; //no move
		
		//------Update-----Base that mario stand on-----------------
							//update for wall,     (I intend to write the code repeat triple for easy to detect bugs)
		assign mario_base_next =  wall_turn_reg & ( mario_x_l <= wall_x_l) && ( mario_x_r >= wall_x_l) && (mario_y_b < wall_y_t + 5 ) ? wall_y_t - 1 
								:wall_turn_reg & ( mario_x_l >= wall_x_l) && ( mario_x_r <= wall_x_r) && (mario_y_b < wall_y_t + 5) ? wall_y_t - 1
								:wall_turn_reg & ( mario_x_l <= wall_x_r) && ( mario_x_r >= wall_x_r) && (mario_y_b < wall_y_t + 5) ? wall_y_t - 1
								:  (~KEY[2]) && Drop_reg == 0 ? mario_base_reg //this code is used to help mario jump at the edge of wall
							//update for pipe1
								:pipe1_turn_reg & ( mario_x_l <= pipe1_x_l) && ( mario_x_r >= pipe1_x_l) && (mario_y_b < pipe1_y_t +5 ) ? pipe1_y_t - 1 
								:pipe1_turn_reg & ( mario_x_l >= pipe1_x_l) && ( mario_x_r <= pipe1_x_r) && (mario_y_b < pipe1_y_t+5) ? pipe1_y_t - 1							
								:pipe1_turn_reg & ( mario_x_l <= pipe1_x_r) && ( mario_x_r >= pipe1_x_r) && (mario_y_b < pipe1_y_t+5 ) ? pipe1_y_t - 1
							//update for hole1	
								: hole1_turn_reg & mario_x_l >= hole1_x_l && mario_x_r <= hole1_x_r ? MAX_Y + mario_hi_size
								
							//general update	
								:  (~KEY[2]) && Drop_reg == 0 ? mario_base_reg							
								: BASE;
		// the highest is always equal GROUND + MAX_JUMP
		assign mario_highest_next = wall_turn_reg && ( mario_x_l <= wall_x_l) && ( mario_x_r >= wall_x_l) && mario_y_t >= wall_y_b + 1 ? (wall_y_b + 1)
									: wall_turn_reg && ( mario_x_l > wall_x_l) && ( mario_x_r < wall_x_r) && mario_y_t >= wall_y_b + 1? (wall_y_b + 1)
									: wall_turn_reg && ( mario_x_l <= wall_x_r) && ( mario_x_r >= wall_x_r) && mario_y_t >= wall_y_b + 1? (wall_y_b + 1)
									: mario_base_reg - max_jump ;
		
		always@*
		  begin
			//update speed if the KEY[3] is pressed
				if(refr_tick & ~KEY[3])  vr_next = 4;
				else vr_next = 2;				
				
			//initial 
				mario_del_jump_next = mario_del_jump_reg;
				mario_del_run_next = mario_del_run_reg;
			
				if(~KEY[1] && ~KEY[0]) //if two button is pressed, he is not moving
					mario_del_run_next = 0; 
				else if(~KEY[1] & mario_x_l >= vr + 5)
					begin
						//update move backward to wall
						if(mario_x_l >= wall_x_r && wall_turn_reg)
							if (mario_x_l <= wall_x_r + 2 & mario_x_l > wall_x_r - 2 & mario_y_t <= wall_y_b & mario_y_t > wall_y_t - mario_hi_size )								
								mario_del_run_next = 0; //mario is stuck		
							else if(mario_x_l <= wall_x_l - vr & mario_x_l >= wall_x_r + 2)						
								 mario_del_run_next = mario_x_r + 1 - wall_x_r; //mario is shifted with small distance					
							else 	
								mario_del_run_next = vr;
						//update move backward for pipe1
						else if(pipe1_turn_reg && mario_x_l <= pipe1_x_r + 2 & mario_x_l > pipe1_x_r - 2 & mario_y_t > pipe1_y_t - mario_hi_size )
								mario_del_run_next = 0 ;
							else if(mario_x_r >= pipe1_x_l - vr & mario_x_r <= pipe1_x_l - 2)						
								mario_del_run_next = mario_x_r + 1 - pipe1_x_r;							
							else 	
								mario_del_run_next = vr;
					end
				else if(~KEY[0]) //moving forward
					begin
						mario_del_run_next = vr;
						//update for pipe1
						if(pipe1_turn_reg && mario_x_r > pipe1_x_l - mario_lo_size - 3)
							if(mario_x_r > pipe1_x_l - 2 & mario_x_r < pipe1_x_l + 2 & mario_y_t > pipe1_y_t - mario_hi_size )
								mario_del_run_next = 0 ;
							else if(mario_x_r >= pipe1_x_l - vr & mario_x_r <= pipe1_x_l - 2)						
								 mario_del_run_next = pipe1_x_l - mario_x_r - 1 ;							
							else 	
								mario_del_run_next = vr;
							//update for wall
						else if(wall_turn_reg && mario_x_r > wall_x_l - mario_lo_size - 3)
							begin
							if (mario_x_r > wall_x_l - 2 & mario_x_r < wall_x_l + 2 & mario_y_t <= wall_y_b & mario_y_t > wall_y_t - mario_hi_size )								
								mario_del_run_next = 0 ;							
							else if(mario_x_r >= wall_x_l - vr & mario_x_r <= wall_x_l - 2)						
								 mario_del_run_next = wall_x_l - mario_x_r - 1 ;							
							else 	
								mario_del_run_next = vr;			
							end	
					end			
				else				
					mario_del_run_next = 0; // vr == velocity run			
					
				//CONTROL JUMP of Mario
				if(mario_y_b > hole1_y_t + 3) state_next = 1; // mario will always drop when he in the hole
				else if(~KEY[2])					
					begin 
						if(mario_y_t <= mario_highest_reg) begin state_next = 1; Drop_next = 1; mario_del_jump_next = vr; end// when he touch the MAX_JUMP_ highest level he will down
						else if(mario_y_t > mario_highest_reg && Drop_reg == 0) begin state_next = 0; Drop_next = 0; mario_del_jump_next = vr; end//up when press the KEY[2] he will jump until touch the MAX_JUMP
						else if(mario_y_b <= mario_base_reg - vr) begin state_next = 1; Drop_next = 1;mario_del_jump_next = vr; end //Shift him up with vr distance
						else if(mario_y_b < mario_base_reg && mario_y_b > mario_base_reg - vr) 	begin state_next = 1; Drop_next = 1; mario_del_jump_next = mario_base_reg - mario_y_b;end ////Shift him down with  small distance
						else  if(mario_y_b == mario_base_reg ) begin state_next = 2 ; Drop_next = 1;mario_del_jump_next = 0; end // he stand to the ground and wait for another press key[2]
					end
				else if(mario_y_b < mario_base_reg)	begin state_next= 1; Drop_next = 1; mario_del_jump_next = vr;end
				else  begin state_next = 2; Drop_next = 0; mario_del_jump_next = 0; end
					
				
			
				
		  end
		
		
		//-------------------------END  MARIO--------------------------------------------------------------------------------------------------
		//Color output
		always@*
			if  (~video_on) 
				graph_rgb = 9'b0;//white		
			else if(mario_red)
				graph_rgb = 9'b010000000;
			else if(mario_blue)
				graph_rgb =9'b100000000;
			else if(mario_yellow)			
				graph_rgb =9'b100100000;
			else if(mario_black)
				graph_rgb=9'b0;
				
			else if (rd_pri_on )//& pri_turn_reg)
				graph_rgb = pri_rgb;
				
			else if(rd_d_on & mst_turn_reg)
				graph_rgb = monster_rgb;
			else if (rd_c_on)
				graph_rgb = c_rgb; 
			else if(rd_wall_on & wall_turn_reg)
				graph_rgb = wall_rgb;	//red
			else if(wall_black & wall_turn_reg)
				graph_rgb= 9'b0;
			else if(rd_p1_on & pipe1_turn_reg)
				graph_rgb = pipe1_rgb;
			else if(hole1_on & hole1_turn_reg)
				graph_rgb = hole1_rgb;
			else if(rd_mus_on & wall_turn_reg)
				graph_rgb = mushroom_rgb;
			else if(rd_goo_on & goo_turn_reg)
				graph_rgb = goo_rgb;
			else if(ground_on)
				graph_rgb = ground_rgb;	 //black
			else if (rd_c1_on)
				graph_rgb = c1_rgb; 
			else 
				graph_rgb = backgroud_rgb; //background
endmodule



//Keyboard driver
module keyboard(reset,clk_kb, data,up,down,left,right,fast,jump);
	input wire clk_kb, data,reset; // H15,J14
	output reg up,down,left,right,fast,jump; // pin led1, led2, led3, led4
	reg[10:0] data_reg;
	reg[3:0] count;
	reg isBreak;
	always@(posedge clk_kb, posedge reset)
		if(reset==1) begin
						data_reg = 0; isBreak=0; count=0;
						up=1;down=1;left=1;right=1;jump=1;fast=1;
					end
		else 
			begin
				if(isBreak) begin //state the buttons is free
							data_reg[count]=data; count= count+1; if(count==11) count=0;
							if(data_reg[8:1]==8'h75 && count ==0) begin up=1; isBreak=0; end // I 
							if(data_reg[8:1]==8'h72 && count ==0) begin down=1; isBreak=0; end // K
							if(data_reg[8:1]==8'h6b && count ==0) begin left=1; isBreak=0; end
							if(data_reg[8:1]==8'h74 && count ==0) begin right=1; isBreak=0; end							
							if(data_reg[8:1]==8'h1a && count ==0) begin fast=1; isBreak=0; end
							if(data_reg[8:1]==8'h22 && count ==0) begin jump=1; isBreak=0; end
							end
				else 	begin //state the buttons is pressed until the break signal occur
							data_reg[count]=data; count= count+1; if(count==11) count=0;
							if(data_reg[8:1]==8'h75 && count ==0) up=0;
							if(data_reg[8:1]==8'h72 && count ==0) down=0;
							if(data_reg[8:1]==8'h6b && count ==0) left=0;
							if(data_reg[8:1]==8'h74 && count ==0) right=0;							
							if(data_reg[8:1]==8'h1a && count ==0) fast=0;
							if(data_reg[8:1]==8'h22 && count ==0) jump=0;
							if(data_reg[8:1]==8'hF0) begin isBreak=1;end //break signal
						end
			end
endmodule



//VGA driver
module vga_sync 
( 
input  wire clk, reset, 
output  wire hsync , vsync , video_on, p_tick, 
output  wire  [9:0] pixel_x, pixel_y 
); 
// constant  declaration 
// VGA 

//0_by_480  sync parameters 
localparam  HD = 640; // horizontal display area 
localparam  HF = 48 ;  // h. front  (left) border 
localparam  HB  = 16  ;  // h. back (right) border 
localparam  HR = 96 ; // h. retrace 
localparam  VD = 480; //  vertical display area 
localparam  VF  = 10;  // v. front  (top) border 
localparam  VB  = 33;  // v. back (bottom)  border 
localparam  VR = 2;  // v. retrace 
// mod_2  counter 
reg mod2_reg; 
wire mod2_next ; 
// sync  counters 
reg  [9:0] h_count_reg, h_count_next; 
reg  [9:0] v_count_reg , v_count_next ; 
// outpzit  buffer 
reg v_sync_reg , h_sync_reg ; 
wire v_sync_next , h_sync_next ; 
// status  signal 
wire h_end , v_end , pixel_tick; 

// body 
// registers 
always @(posedge clk , posedge reset) 
if  (reset) 
	 begin 
	mod2_reg <=  1'b0; 
	v_count_reg <= 0; 
	h_count_reg <= 0; 
	v_sync_reg <= 1'b0; 
	h_sync_reg <=  1'b0; 
	end 
	else 
	begin 
	mod2_reg <= mod2_next ; 
	v_count_reg <= v_count_next; 
	h_count_reg <= h_count_next; 
	v_sync_reg <= v_sync_next ; 
	h_sync_reg <= h_sync_next ; 
	end 
// mod_2  circuit to  generate 25 MHz enable  tick 
assign mod2_next = ~mod2_reg; 
assign pixel_tick = mod2_reg; 
// status  signals 
// end of horizontal counter (799) 
assign h_end = (h_count_reg == (HD+HF+HB+HR-1)) ; 
// end of vertical counter  (524) 
assign v_end =  (v_count_reg == (VD+VF+VB+VR-1)) ; 
// next_state  logic  of mod_800  horizontal sync  counter 
always @* 
	if  (pixel_tick)  // 25 MHz pulse 
	if  (h_end) 
	h_count_next = 0; 
	else 
	h_count_next = h_count_reg + 1; 
	else 
	h_count_next = h_count_reg; 
// next_state  logic  of mod_525  vertical sync  counter 
always @* 
	if  (pixel_tick &&  h_end) 
	if  (v_end) 
	v_count_next = 0; 
	else 
	v_count_next = v_count_reg +  1; 
	else 
	v_count_next = v_count_reg; 
// horizontal and  vertical sync,  buffered  to avoid glitch 
// h_svnc_next asserted between 656 and  751 
assign h_sync_next =  (h_count_reg>=(HD+HB)  && h_count_reg<=(HD+HB+HR-1)); 
 //  vh_sync_next asserted between 490  and  491 
assign v_sync_next =  (v_count_reg>=(VD+VB)  && v_count_reg<=(VD+VB+VR-1)); 
// video on/off 
 assign video_on =  (h_count_reg < HD) && (v_count_reg < VD); 
 //assign video_on =  1;
// output 
assign hsync = h_sync_reg;
assign vsync = v_sync_reg; 
 assign pixel_x = h_count_reg; 
assign pixel_y = v_count_reg; 
assign p_tick = pixel_tick; 

endmodule 
/*

*/